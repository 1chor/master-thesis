`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
i6R1spORcwyN1lmmfEySpXbgci00dvotzo2XDqM/7zBHdAnoqwRS1iVz/htxeRIiyMIqQXT6Bl4q
gJYbhcOedw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QlagXI5Cue5NzPU01n3ZmKVrVpMlBDK3ZGjdn3MsSGa7X58hfO4Bby9RBhEFLBNzAOVgdWgxCZ6H
1MH/gqOAxM+4hLqjOn/zyraS1qx0tLTyW2M6F6Qk6UBfbqdo5qrHBWVx+BtA8pUU094yB/YCUs0+
uTmPICZlcVO+3ndtoa0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K7xYi1L6RbJsblSFAIIK2nlxpnIVAg6vY6xNW/3tC9t6bYrRMn81WCHyI/nu8aDBz+5s1FvR3yoz
Nfzw7O61G1fvw4lj/CW2Rf+bZAQFFNMO7K7kPJsNsXBQN690Cj+jSSTXEWn3w31S+UNg6axE9bkG
sQ6Ryo4UOKayB1ycA08E66T2KkWO29sI9zDSxznEiGbbSzsFb7roNaSliVZDbVZSWCQKGQfRW3Pz
YUUocNuJR3K/7CEC9DfGtN5d0SCMleCV+4hmshc/VLhJFudwzhw5CefQiCRkj6UZ0KfmXN4pTBKF
x1hj6WyftkfalWR6G1Of9V2RmreVo/tKe4hJMg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EJo1FlKUEKAxs3UAtHLfZRNNLFxICzGCyr84gCuLih9ZNbtsAkli1gHwzgvY8UfVQgSkJMIpfSxI
CB0MwH7XxaYQl0O+NrBdwBc958pp+XLHqouc2YomENWCgb1YRKXLXC5i2MXyNxPZSFVGn+oEOWG2
UrC4eTW3C/eY/4PYvI24Jc1v1YZTnKU2Pmr9jGHZDGfiD+NJxi8YyDHY1ks+9UE8s0VtWmSNd3ox
UH9c22qaVhsoLqpeXb5Bsu5f/Jl4E7beFopZ5b8FCq6kXh7aV7UHS672vLr0kYJ0tVYIrvtxMXVJ
bt657seLD7kOvgUGuJNDwUImG1jT/3pIn0zVfw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
meOtD6iosVb2EMriI/7eiqpFPX2v4S/3wVI5YoIZ+q/y4KN31hHFdyaiLfUvRbeyh310iYvAE5Yj
n1p0ltmLD/GsCYp4qbMm1cwJ7gg5TqIAWpVDoZiSrYW+bczdqxq+nw96J2IADOBQqTvDvRVt9l3P
EB+PLNzwRXxbS91Ru+vpp18s/DaHzH7D/Kq3FQ+0atF2ehI5W3KKeNbjS5c2VoMREsEf0w6jbk48
54QS0NmTMzg9PkeaYqQz6OdgqYDKj8VWOTRzycnDDyftSbthoRHSeVxd54LtD0sjvv4MXLjqc/h2
+dv08O92LZA8EpwL0qIvyi9fqYKbY0MQZGPdxQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WDEzRuSWJ4Bgf9QwQAu4iuMat4z91QMpm7UE8/JIbewkblGJ/cBiG3DIqmd7HXGp53OFnPdiP5ZK
Osh75v46iQfkU/v/T+bK9Iuj4ZiDC7WZZblM5A2QPw/vlUcAi7Za0j4liOEEXO9qDNVeK8FdIHLE
oAEogzQMM3/6WJF6H8Q=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j6V1+x7/T1uLedHK6l0KiBESl2DV5NMeqGR4jnqzk4hCiChQdleGsrObJOnoACak3PMlQQmuc35v
XjhfHuhkIhXoXM3Li+kv1kljBEId4MnCcHyIeglektFw5kDR/arXjaFOuUCbsPJXwgTOXdjUBJYl
P0mOx9AFWdOHxHDzMPhdWnuLnSBjK+UKgKAIvCLRez3+QwRhDfA4NyDZjcQUcVRWAUB3KHDO370m
2bLG3h4mNhyfG44GLT4lExBhaVwH0be/KFouL6xEWvvQNzn6+SdwLrOfzXMDwX36A/vnVXMF/I86
Yem1uvf2b97oO8kFf0+u8V3idHN4eiPmVV2eWg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 665856)
`protect data_block
RskW2MktgoSh1LHXIvkOWpx7o8t4osGtR/LERqYpeeuaDBEv3QEnXqYrRXvxKgcy7/mhpm8s9TZs
oCJmoUudL1x1o8vsGiZYdgRnX8b0vznXF+bs5mhNPNA0bTWD0dqAGHo6GEon2YSsYZ+fT0LQSUKK
geQwJ0oLtnRuC5yojVN7kGpjGXKZs3INi0yfWQSclN7pEZY9dAdQFiLwgwlg/A2TgDodmohv9Gt9
yYX+OtwyhbRORJv+U5utQMthk6zOVA/vTX7eAt1e160IBwLXYyqSgBMpMptp2Sy/AuT5hLCoKY8C
h2c8a3H6H5BDz9ajP+6OmIBSxLtBZkxiwLBrl+AqYoxQ/sE6/6pGw+9TjW644Yk5JbT4lYVWFk5Y
8VJpWzRqkoDyF5yKSmgGxcdiz8wW9Mc+4RtNfEWCcZWWjPPNC5GeU/qcGG+OQ1aBdwRgwJJiBfpj
DeSaOajJjVHvcmPtKpDaPaNKv4ExVWLbBPO/ybVDJG66QeUJugGS7p77bqHxSjSoUt7So1+vBQ4G
tP1OnB9AS/iePA1F7aqs5luAxITauHHne2kdK6xZ09N/x1cx31eXlpXb+/W2zunoEB52konv1p76
zvnp843a74bHAtxKAzPsytXJekjFwLlAjugAAe7G7MNrZoKRxr/sNHQasRz0Yy02g1HsbzhT9Nc3
L6xnr4HZAWyHdJ6vF8atzNsVLHOvCu+xa4ccSCaz7XfHWcdJ7/z4C19u/0UtmchXzdIfM5OYj4vq
BKWl4/iC04twg5fis5c0+eXUrikBpkRTiLOX8X9zq9fzyLkcZgSn6WGbAF6ao/dDNQFt2Aopn8cv
0RDsSCayciMpGHeh4Qu3aHxSGkvoTzklQXYU3e/4haLVK7NihnKVMw79NNIC/oYzDAVh7GiwIOTO
8xmnMnaUcs/lvOL7PYWjVi/7ATydys6w5uHEPcP2RzM+qPyFjTWt5I+Ss24un6MKF2XMF4cs4j6E
QCtAfdufu33HPgCoR6Uyxjjq7n5+NcGiDfZxPH43DC68rbRnOOW94cSVkFlmS96Hymx12cdImTCu
H4vrXVIXiINIb0g5vF7zMZv9QYVrN+fAEfLnjmwF3tUOy/piNeJ7DWTfSa8tvE0f+lRvTUG9Pmg2
WbPV7bzaIIXy3uh3DLs7+MAeHCRVriqBjRD1wxS5oPnlDzglFcoM7f6jpr1W14tUXmQINV5gG/3u
l5DwVV3/iGhlHBmwhwd9siIvEfIneVBWHfjGMBc45aO9joZKHJ5SJ98cT+NyaDGmkSXVLRqv5UXu
tx9mUzw2KR8UL/5JZJ1O2koA7uMNUf479WVBKe0irMU1TwIL+xfPCW6nfXFlyAcHxl2SV2MtyZzF
4/OXyAaIj6e1rSqTMoBPU6KL0afRXx2EiU2jdaffY7eL3zlAzKrx1bXRqxezWJdxE3tXOYCHiQeV
nCAeWz4Nj/AeO/1uVm8dliwkphpJj5gV6DY0noJFfHkVOfKIZnCwZY0668IReKlHnpJbv6KF5Dtq
4zGpqC+KT9hfICYlg/hQ+2FdqfPDIhb0wNScrlv2B30zD031rR6PiLDZGqVKK0JvqooniXJ1A+TV
Ile/+3ll2LSu4oSqjpVJp7GvLPyJgpL6tngi3rXaN8FRE9E0yIGW6rWX4v6Qr3w+DP+QbkLISPn8
M1/+ctm2zRizGU1tCD2iwK96mfz0IqWTrM3wDCIWIUQ/Qs+NznqRuq3EsZcelmPBQvzX8ytCNJT2
7tWsRsg2a/Fo2j7f5G0f4heOIPE4ElKmc5WAq6hdvOD84tht/M55xnK9udt1CtbOECId8ZJH0IpT
vpJTNTlV9mjFaebwCjJ1nMHjf4uDLPppefqgWhkaHmg3ci3gEmcsER9R9OXGUCgkQ/Tcc8cax3NR
5PynUS/29khzfbJ1+MjIAtDOysfyKOzjIZl3v8Kjk+JcqPh8hiEUXJOFTKi9xI8QChpNHZjkCzK2
kcnOJjKkJpPUzmw6VnqrWvTyMrhjUm4qP/Rem2XEWDU5Edd2i5S4APQBlLGPDioikoRs3yRxrO5M
ey4CO26NNvKQLW5oPT3ItarZDblU0L5b+wORIRoSgkt5RTnOGJ0LH02pLLOjbhpug9dFJcDoriuf
ZG5LLDVOwdbfbWItJNwP+tnRJfujLToDODp5sNGfLtKnL7T7i85eDG+VJbOpq8Zaq4lFloOugN4k
v5ehXf2BEKDJEZtRB81P7yG9kSdeIHjGBklaZHTyZ1rfuPh9vuapMeLXKBkqddFyfhNOG93BPp1A
9h2yvAYX0QUaMVQwvtYUc/BleoS4j21QXnzH+kVFxCO/Uhj2I5uvC+jJPolI6qeYukbAdTn1ZlB0
8PGZnUlJQSjN5eHSjb3lr66d/9VBWB/mD1TWOLNXh+0JHya6obbp1/b6m+gzz+ijY0kgmB8U3kDa
9ZiTmttaZXUiSCCpQOfjKnLsmx30V9OsfDPFYJlrbu0gh+POUBQjWsn/HeB5bY581gVJVJ3b9NzY
RvHk4+IRN9AkAHuXY0AQH+uUFULXxbLHyoPMECdG9Wr1BEWz1luBcriAV4akn59lVV5bHGBat9Vr
x8V7I8YbJCtplKkAvN4cII6RTIj07uhLWmKqgBtm8GU3v1o+XEdJNEJxBt8Ci+OBHN7icCtqAT9Q
kvvBJEqxnfJ0MXMf0aCYNhvK8uoFgLw+zRNYqMHPB6CUZe1BzD8ywGWsABv7lPAvXnXMunnWtn+o
rBFRqKtGAkmAK5roY2QANQXFLOwAxMpcv2soaKzOhkIfyUfIZc4FrYEJzF8RnI5ow9Kdr4UnTT9j
/4inPoPk2KIgKe1BeQCszdRRr4nqtwLWp23W1X/Mub9rd8W5d/NWleMh1AqsVLZoNsUb+Fiz8pop
8d1kQhHDW8QjFd6RA+sQGZODpkdkD2CDLiwsDvc20/CD7k8tHlUecewo2E2UG+hXDivMvn9AXhC4
qZ/T05ykgwUkCPsYk6p/NdTTvrj6nfqge6aPzfisepkbA1JVFnGK6QcJMWR9NSn7ifG4vj4NJuuj
LKtmiWX10+t8GwqWKXp+CrZTmptZEXvcjNT63bmMsFTbKzHVmCEELBCi7/fsmOjjn4pnwpiE3/Wq
mHp9cngjZssyakfjYvnqOUkXgFpYpA5cwg22sSa3tQQ9r3a4vzmnMg/72Gj1zLGo32b5X11u1Ipa
z91c6iYO9/RK3z42uKyJfzYwdwnV394TJoc43/aPW1EyLgyu1dl7XuiFUqQ3/H1QRdnHTJpWbG6g
N1K0cDnzw9mU6VKZ2ZK/8uz219B2qaHtL/C+4RsFXKDq8lNAR5HL90xGC0aKqePTB2JykP+9xvdb
Xg6MjXdRhPWrOgAIIrmT94RzJ5DDOgcquuR/KCQqoLcCQlU3U5cGIfIjvs8xRxDlVTxkHHg1se+j
Im9Wx/CoLgdjV1iBAARHto5nPfaQz18fp9kLPKoxgn7L3uolrX7eUIEX4s4I34OIBuW9zcR9SWxE
Tw6D6xYF81J8mvDwtL2hO26EFsD0DbmIHVitUgG/VOgnFb2kYi+5SvjtdVsMSxL/ce47Tl6V77HN
4lVux9nexGIhBK3Ot8+z4J9N43+z5srcrkP4PORwu9NbcZDPpAVLGyMFqhso3vcQ2jDLR/a8ryGQ
dkL0g8ayZ4dwNNd2OfT2rE96yPA9qpjaXNh5Bd6obFVqW3VBDMOquKtsZH5xyPPNwRpC2FmqCMfc
1rL2jI3bZzPwHyySfaWop/06kF+u+0L3nXyysAioT699vM7VLjXhwMbMJmM/11L7RXTks3uaJgoP
fGSD9n3BtL5lIuqXyZWEjmdVYCrvUFMiFHRLdQ+qaVgv/L2C85ndUX/amraaxHnEuRgZht0GAJuv
9/PTFjitACFLyYOPaawWeUsDb4dEymSF9bxxxU2vIoYLv9bMOsGvYU1kl5rrg6CoXQX00B+Ji23J
vKY5aUEdgSE7OYTmMh3EFpdljMXYjHeQy75OYQig+udlogailcK4rmSx8TrZkZbdBOliKMtKCJrf
jbP/m4swdUhq7bggxyOI/2Jxax0iV8GR3nap/dr+IQoHQJNFughGHunKQEnyKk8Wkk3ylUS5y6iK
76ECGElfK+z7SQWyfN+imk6E0aVAhKhZNQ4hc0pieTJnOOsmmJVNTtiJeULetfgsHe/dWmDNLqUL
koMe9genlNEZSbGWb2eZnNSyQeguuSZfNxwzCAYH9Z43B3FqzJyMRZrtkIbj5Aq6haMQdXkmmpn/
04debajjvnwkHMocgy+Js9ZQPEGekn5K1C2KtJaHNM2aqHK7L4GDTOrB7V9T9evaRdCIxmJ62ype
zJQLt29beY9ASR8K2UNib1h5iVGV1p6/NW3VvtVAZhAknwtbnR5zG2OhzLAmaNA+G/ks8zvGsdIl
vkMWoHLIpUR7aLByl4cRQ4WYwmR5NQ3N27T4Yd2x88WYyZ8T4Ban3Wltn6Mj7rPnkA/LlbCFuQ7p
ZXl99RClFKBoAx/dS9dC7oMUgFr+fGlRN1xGnc3ZfUYUMlEb1QMtgD8zX2KkMlZ1G9wQWWzOrlsf
9uQ31FJMPKC9XwR9mx8vaAnBBzfOTDNEKAAzQevEfi6vpEXl8oVSbmrsU55y7BT7uqQS0mudS6Hv
Gp3LPiEYsNIkSmXfDJfkZWWAgmbTRQUHS1tcPrgOAvQPjqSLL33jmyHE+oE4CMjKl4eJhMBUg0Xs
zwbOQbAK9ot5zwJvgcuXLRdfJC66rxqOSR7aJidICQU5TbjjQkYqDazfIJQqzNjpusApWIEWY+84
xXRpjXWeD6Nf5tUm3+NYOUvILZyktM9z/z7EL3QcEsL3P5ggqiQ9cLLgKp8GvhM0e0wIEuva8jMF
/sCqO1JNmqjStMHImr8olgIOMCfGj6W6Ujt2jevb3/773Ly1d3AsBQm20ebbftY/2Vq9/avXGH6j
nZWWAZk9BVqVqbpeLMWiukEvLlXLuOf9qAoQ0KrqNaf5CsJE37bGX/z20Xo4OTEQj9Y7bXN+8ys9
Nwx8Jnv8X8ELNs+Y2NtirrxTgP55CaMcbeTm/dk692pTmgsqX84QsEOlhEwzKQDwe7Rh4FvRIYg9
OvoH0vEpED65baY8cAxHfLOFAPg3LyhhyAViNkXPToy0uodTuhIL8H4IasK9AmzwavbaPSvKRG6l
IdiJWSxaJZnXSYUNkxNDkBRsskPfygNr4/mdEtPa5LbyE3Dvu0ZzVrRdq7kpaCQmKJQSvtsxrnaz
Q5zjQh7bGmTNfFM+jCM3ANjLi/0FU/CWis0W1D3of9TpJsM9jzABTtUEEwMAMFK5kfRAK38f/UGF
OIFgsMV6ULgTPC3cVnykCfghktd6JWS5y2KdPa6/WBvTa0dEhW0ktkwdmMLcdwHMftABTmLbOBih
QVAjK8+swZ/64Ncz0wT1COFaM8xGiT7+d9GSl8ioOwhr0kBZPOwyCmrEVbQvtY0VGFaf8kUbmFIO
95qBsY2RUxV1j/GE2AYjBYm4NbIGimKLOYLJqD0NDgRaYV45DX2prjTOO11F+zlTZPtVh/lZXjAg
F4DOAFVuCbtltvdxtPW4rQXBIZ66lvzyYM7lrWOeDz6chrNfixF6fSL8OYP9USeT4HDER6aCfmov
8uS6iHKv89gPpgx4Avgb3QovDT3OZcFEdU6f3yzGYIg+7CvOpe1gllz9G9zh+D3cgRvOWge0VqGb
tw7EC2o8W2inaKZ5pvYzEGeyruilyViNdoOqt33sQo/4tV9eSkVr+S2sev53y+ZpOazHa+wwB2nd
foC5MznZbddPM8NLIfcGlqPIEKb+OZlrhZP5inqmgvH8rKizgv9JwUUfYXupMzuRt50Rl16coS+6
ckjBT9nTLGELcdVwM27mf6f/L6WIgR/b+EyWSkPxpSXieel8HUsRfA9p8uEXIsXm1FSsEP0eg3fZ
fuKqZsm6hnJvThN8LiJXFWglgavyzJOJ3awimjfknSElQO4mZ8xfKDvL9dKf6QyAUV3x4A4R0Kms
yJ/TuhGZH6llYQUFox2Sek1TndO5TMRS3TGkeN1RzksUah+Oj5gj3o2YyhLnO/yKcIXefFA1a5Xo
qGwelvmaBV+ZkvejckE9UrKDdMJ5cCMrFjVvxFPY0enFhxNK60ebZbsSz3V+BHXi1FmOSGSBFroF
O6KU0PVC+PkZ+o7hHrNfOC3hzW6ibiBUu0wC6u+GOaMNHTVH7ZZbq4lAI8GKysaWfiRettSyQQVv
Mu05k9ezd7JKLKAUhtGl0eAfrIYDtxu3TqlmRREXKQyO5kQuU80kwRbY/O21fZEGc0QpcaoEhc7w
Am6VGLsEdAVmcLZJXj08LH/0WfZvsJz4uSVUw751cagTM240ERJbwpuUGfDmOQXKczQiS3yqKg4m
jHcTo409X0IFAlDKSIQ8fnkvUDwDpMCQUcN8abMiLjgYNSKgpbf9/GeoqKTAFtPaJWzakX8wzbT9
4Kk4nVYURIcsm+cTu4EMYeG3gA7A4eVrwlLSE7wHba+mt0C7ried4tRKev/ELfKHcUBvHKKB4kta
mVssDXn6HyBzFdTKBQNlM0ijDJDDhxSuMWK169JtTDdsUkaqjQ6psQTYEBbqqlG28nql+5fahfYU
PU+wNm2B2OwMfXpaE47hyeKkt1iG+kQe7WRmEjfe6JvYlo4A04Sk6Y9r0Ohl3GIuvDPA+5saamvu
fl5e5kyyIRz9NClo/qwVGXXVGIUMhlgJEpk3v0amhH6vC8vWt62Z3BQMj/1C+3Ykauk69XwBuzYx
JsTc876y4E0BbJm0P0Fp2UdPi1eTiaCQXDL8zMY23HWlKNIR07PBmRlIwWgFmh9v4Wy+D8lRuJLb
HjlcoWRDlhh2H9tlUc41T5rX4zkl+Puvd09OQvGnTN8EKJejUT4loppXz6xufAV2H1IOYgo+VvCD
Aty2XAMrJhhumXm0N6zsgw8xuM4YqTXi7mdZTMUzQUu+bPYjKCgRUyTWkKBqGRIKSGhbiFXDX6qN
aVcHnBty3Dlq/pvCuwwqiVeZ2P7mzsu6UiqfNJLYaLGeR+ZJDB6OQz+kexT2H0HS74AfPIPlgsCC
1fIXGdXzjzBMjs+aC5qGo/Wec3/04UUXE4c8uUjr2WRAphbGcz9DXEXEE0qGhC/9wt8clNndPGMe
bRWxWTfQ6LWN5C2FQUO5Lxy0Fh9L80QENDznuAg8rVvmIxlIa4N3+YHlgT7GICoakhyK2K9JTqgr
nSyjxOG46/7wIyK4dIz0gSYo2GTfh67FsDkgLjMpPoe0qww1q/w4LqJ5a+4rMOEH+4nGPBL/BI9C
IkORXwMxraa5aNLHBQ2lDo3kYLeWihXjp29L0pzxVtKO2HMIzzCj3McXeiRBuISuqxOfUO+KM2Q8
mCC2v5nFxceeL+4NwffvtVHQ5KB9gLKY5kj/AaULgKHZtluL0R3iIqjM9Zb2RffjvO+LF0JNNeuv
Zjjoio2LbrUTDA8quPc1xXDMAxiCxhYpGHFuPd0A2ZkEYBt+epdfoLnvhTBKcWLsocBvi2XdXEtv
Zcp4/k6KYsQGjSJ1qk5NhO4iRl3nY3pU8BFfc+yjGEd4hU7XPsm4KkPLrvJPsmvljtOt8pj5hUdB
4TB7tGH3fmYKNcwnU5QHCWlnY36EnzkQ4SrKCUktzNNWXdblroOuFaVIAT7NMHngINrliMPlPun1
rxXG1mD8GuezjM1iLDBxMPvrrkhdU0hcCApOYA4uiK9lKLm+s8JBU22Ufk9OzwCpEHRFalY9btOd
ezpXQy57GCjbNFuf7XDgNmR02AQezj6UFbxFdreD0drTNWMI6f8s/Zyi69eWIePCRZCEjIUlt48C
swoW22AbzkukDPODQvVqWD8EuoN6kwWe2j4eB1HgutKK3HKpNBB1sXm+Fn8a62O2YXQOCYV9JReu
nRC6YuPg/kboCC2UG2AO2TTD9TRmM1ekxN0nZtRiIZjCuJ3OOVr0PGiNqEQ2pJ1q0avh6+746haP
6RDUMWrA/ZbxKkjHGXsG3ag1pOEUQcWatVz4EJ2jvqfWRxi9MKPG6rkcnRf/mmaKpKkmZeQpPzxv
Z3JZYDPw7ebEs8KaXbStk3zzY/rxDQAUxznt28S/vblrv2+1rBanurkO/ft/XzlykD1ep9f/dBlE
9ePsnyFz50ybnz147WJHdrP6b5wuT1waUvEPjcVZUYYrqmKLjV9E3A6ZHIFWlJQIR4CpoQHRENhw
isBjgc3D7l+ExYeRUMn7AEtVtoKKyZKE+FnEO1TfC5VsFYirMl7ZbTYfLXuo2ajxfJ3q6iHuPhfO
wFj2KXOxKWqJ41FuyFDJdSEKqXZOYuJF6UtloOmpQ3KZrSXSijGhjbrnBP1KxCT2KaNBRqdJHMXc
ld8cR1AsFqqLlAfSu9BtxMLR1iSC/nXLqAcRtmetYY7WMap/CTbYJsoTBnV7qSoyM4hqAhzWc/UF
vAznTS3c0zbMJOAHGlwxtjIAvDxAOUGLpU/ZT4hrLDb6JVTpvfvSjyS+f+sydpsi+pNwNjJK6vkv
rMYLxR34oIJ2b4RoviYF1BMcrQ0AHmYGXXeE67iUXdBdDZ9KHBWOse/zf1KqYMNtQJQZigVKCxGp
u5kyBn8Rh1vh+7bynBVUY6umdvMe0JAEhzDvV1GsE6kye6q/KoSIiruNWe7q1/aQ9cFFqfIhlgyV
bfktV8vg9zzaAVabL78UuYgZxfzoMEa5lwWG7bF4rM2Rx5Dmk5ZBKT5wv4AtZf3bMSSVsq7e1/L0
P6gCsbpOi/1JIRYr+cMfvzYsv8iwwrL3ucYmW55m7dPjnWFYHc/hSFVnt4mzIoAmJ5zuPSVE9Kas
vSLL4bC9C+IKqVcs2CsMOf+mpCr1jTWraObYvsC5VU14d9LiUKnN2cV1CfnKhegGA2DPR2wW4rTj
vUMb4oVxOo9Ad+WUx8wKqz1M6dBZKJVxigKcg/pE0T/ifVfm+enFE1Kb3QVYA/yIjQU+Gsxyqnjw
KWTaXr9wtM7RXcFgzSoEb6p6GtJ5/234TGerQJKsAQ4EpsCnuOKzeObMEv0rvrTU+ryyEtXT9H/y
GVXufWEG3g2nVUQklEhnTUVtupep+eCwFh94ZmZT4wZOYhcntDD5u25gbKIEmWaZUUlBLpIRDW0Q
uDunBTzAPoVCDMvsWkDOoftgVOlaUoQgaE9mNEoBfyxd2zow7aeVMfmRLMTvYNNIZ2WZW6xxIbgs
/oUhXqPt37Zp7J6wnwJfroQ1xg/rb1f820EPn6TyqzjRNbvjK/tlJPEMHrhsDxqz+wDu92sON9Kd
jZoaJ89IjO1fioiUt/aWk6WFetD6nE+T2amrq+IqxuVUhMCXfF0SreAmSBSnZJIpFX4wRbD9Xa8f
W+KN6EpwQy+AL0v5nFsF6zLPhoFfIaiwz8sVtE1KtlErC3Sks4BcTYr9oRaNtwuprx6aRof2oL9x
xMYV/dguvqVYhZba28T9J1s0IQgaJ7xmqp1nunsqXhoaXgSCg2IcST8GRj4J3TQhog07HaKic1EU
XBvQe4VqVncKsCGcoqMGlq9TO+WO035GR2Rhep4/yEbGXnJ63mDFSyGLm1NazxIl+3ifctRNm2mL
t4NLvdyEIP/8xwZSC665nb0ppnZwfYRhd07TnZejIae+mlOoL6iZi1JBgzjEDEZvroLyQi37sSgP
6VykeOh01vEt+H+K6CrQB3bhea4lndjLF8zaPekE3L4b/4ikvMlU4FC0P3HcUF5pGo5fAmTIsgrA
pX7VNJG9MIcP9nB4itM10tlrxYd16BQAZGdOlWM10xO87NXP+dm8Ct3XbfQhERNeh7kbIrfK/AVS
hmBhIsMosjP8kA2AxVsuaufuGSkqsFC++HmXX26LD2Oj91LY8WnbONIZP087LvuADcw5rqWeaasp
L37j7tHMShruUl/94NBWHZqfben1/iGeEBdiQT949yQ1z7B64zthdlMz2CiuJ2a1UhHNDw/x1v9X
9dAPpb/oHs1koasp1HVLQaB1aGYeMh6Of4ydHu0Y/tGk5IwXmcc2jIxrsBJgWws3lJYxPdv8viHn
qRKmTYqXEkFSdECTxbL7FErq0xbpPdjaUw/lZ7VfvM73YsURyZVmKtoRXiwlovUqNoSRClwXFgQn
cSpCOcxWNr3VIT7LMQWR4gRf2oUnkUSa6WIQi5ZCsFB/wQOfPUF5rIuH/MWFBclRn+F0jBAUC6vM
qzzVVx/DSIfDl1wPldFTBnbcAA5Sgd132bt2x3Rpm14TP0T51gjRk+KBFm0Hjc2cOfG9++Nnf+bi
lAXav8tHV/DWQQMuXFEaDo9mIZM3vjBEOXkTwXEkYG4Ej9agv1RICziegpMDm3vzwpkFjOwTZItK
8G3jHMOOlbiq5a0rLv+CEJnKgcQDzvdSOPwQMxdVEAdrEEkGF/0rkA0ChTXlig9BJoSqoC5FZOYE
q9jJY59wXTblLBckeCF1b+tIHUVR+kXLcAkR+Ex6skqgaEaYZkVmkDIwvZCOs5HAlHl6T494hySw
L/he/MJJtP9Ge9n9GJZINDZHjdHspz+2t1UMsZMxRd62EkELJCAhILtY5Pp67pEtlpH1IF0L5Z2+
Z3CVhiu4x6fAaeD+jL3RyUNfv4EX1hb+PHE3AsJ7uCcCx5Zh4A+sNw1RrovRlYBYLwPvFuTlSEfV
xkr/dORTpzKV9AX3mk3KnitUQQAJTgG2+BrDsz+KGGNy0142e13RkckcVHQF+xQ7oRUXUJlsKa+c
6Wz98NTfc15wiah/e3yNDNSlNPoTN5kvJ4xacmGTUp998+j4HKuFmewxoStuGAk2J7XFWEUvBTo1
LXe6ndCq5S/dK4Rcp2xSFIPNS5DVJIMG9Jhs8R9BgNgStG9lL1UNjbeHKwQai2BvlQTD5/LhyVwu
b3v6ZHL6LMeQH8S0iObf5ozbJ3q2SnRTcxzetgZ0OQpF4EXWS9V+noJ5sIO5IqFnVhrALwn6GXh5
CTYwSa4ooXMfvul7DwV/65FtrhChlo672YIbyVoE+zet7DiZ8pKj6FT7lIYQpOicWFn4EK29ROZR
XiC3GyeRknAMriFdvvJ6esoX0Tj9+k7XkpxT5lHLO32BEj4qqkAyvhEOvZONJ+mJ1I7cb3QC/J6C
zLGnS/xKYkRWu5k5ksubBhmznl3Nyc7qWGlPxtyuh/U20tpd8SzZrRDVykVjJlOzafYFtFW7n2M9
rAhTnkbpJss603CbQeGwyik56XpA2NJue85gz0GWbWHcwixkw1K6uk7TsHa5KuZvJ09jCeMA3g4c
o9S/5WIXDgTYRGw9CgsqvNkiIoRr81wZrWClqFA259SzZKkfG8jdIbr4gQ1UYNnp+8nZ9i2dHZ8q
ZLViWJMtLUNHtOSZRHtokecg8U6Jw+RQwa9GUtjQFJE/fpvrSBg1/4dPw8QJR2vnAGLkr3bauI01
hh+VXMQcALF7nYwolnT3bhu/G4tkiRzuO5D9UBxW+SRf6rbA7f5Z3f324AnIUWCII4xhkmYMkUFA
X4/0S012pcBKkC1oZX/Bp/T0i6IgkwQ0nN2ztCWNUZMlOMw4oWWFhauDU2a2IebYsMSL9O76rlZb
1CeyYDhQXozbykZl9aTi/kZ/Irycu6FkLpgdeuSfkn/AZznvw7hCIUPR2Z7SeJ80MVNe3F8zsa1D
6/n4aPrVDcog09JzV1ndzUlXM33zhYzmA1Pvh3ljztsVUz4g/4qyfF1RMTZ+8vCdQ1Brv6utQHop
xiviqXZbF0Ym8ri3eoBVHO0beVe+8WqNm2A8WcB5zsVM4Ai0zbazpZHNpVSs/tykxk5DimdiBUrE
78+bEfeapw0+CIQ2Tl5hFcrBMKbYdBGeI3yXTObulHdilUp6CF4/5eyPDNndDiVMnIHYKDi5MAnA
7pJnvOILXGJp/4kgeYV4m2hla1U01C5zw9FsXph3Xc0Xh1Jt3oc5SxHu8W/km4VZN83y22XADW6J
eDdqz7rDByBCmO1NHHisCmVcVH3dZ9NWlVE3kZE+MKb14TODmJ561CdL9O929HsmgrexfahR0yTG
NDOp5SR0D3i0iSO2NY4h923IMicfYotgK6C4o7hTKgZqXF67oU4RYtpMsw4rnRUdBjkTwruB7jZF
9nbxk+4KVuA16EToqwIIkv+z7SW7Ll5k9xXFduwHraZJwKQcLCpqbxYD5wUR4vNmA8oWFU38bDDo
7nMsLG2pZSN9pxJ3rBaACxEgZafr0X5rzPnOcte5+mSkM27/pDeuT/ygACXhEJYSKFMPyBC1OBzu
KhuiXFq/3bnAQ1erHkc/cVnk7ih8Ao/jPF5uo2hf1bGtvJFfTMOOS/OwH6gxZYzPF4fYYEeMK4+F
NRlwjAv1Ixc0fRvRX5LuJpotmWr2nkHeTgecG3ZRmRJkm4zSnECHFRhlkY4WriGdlM6075LajXIk
uya1Sja3Tc0qoVvIvQVHFiP6SbOkRXsOhiepFRlAa5buHrIy3cZEBS9DpiqPauBt7ebfWD6+IKbw
pB3K+AjFrzq4eiszmV27OxhVATNyKgVsoHVhaAkqI/IsImR6cPar18IxZjZD23EG1ceSm4/9a7+8
UWdoFNaAhVMpiUR6yBT00OucFh+ufnXAEfHfsbmJDZEcDW+vmIhJqWNiLXNSGrYPs7f+XMTkTZD3
TyP1AToLOHF19oqgmV6a/JKf8pFKYhOB7z010+1aS3H17BOo3KEAOf8IPFdDD8n93ScwRcP7tmty
rmst1jObLZCRzGt8QV987IqciV5cE5FngD/dgqXdP2Kz65dw55g+UlX905BlNuVTjfeXi+FTY2t/
T8fEziuLeQWJ6HeB/4rVDrjVjiQ7m9GLivynky1CWCTL9dCQa3InzozKLJPNw0RJB6hiDKf9Pus6
6VwyvJ7Ygox3c/fO9z63RkDJaiGOMBAcPwsMVHZFPk1Q0rHWULTCm3cLhKS1n9IPXOlsnEjQ8a4q
gXsVwCsWKrdOmmkXCECmVjR6MLgqw7bxHnt5StbIoNuQR6rc6HEpfmyvuMpoJ2+DMRNHxfLKMLR2
IKkEQJeGIQG0zydcxa/NLoFdT/RTXvMq2A7Abu1zjC2YjeTj5lDThoEDFh8oGpnCDf7I9HYIxtvi
oRQNekE2j7e7DS2QsbiI/wZ7ltSqdG360rcRwOvvEAzVZB5614amPQnyJzeyWvOe6arS8qayQAS+
Imy94qRTiBV1d1grvpzaeoUBC+YRSo+/uDzKx7ADGdzYbvXSF4yoC7IFo7Y/Wlw6ps+GjfDJxwoY
S+Bt2fAm+8eCKMLueZarRrcmNTf7zRCFUOx8S2bpq0Vcj6QSW62BYhyEEBCR9cO6A1rtVQ2ggMYk
nh6TswjRsY1Q3AtW1EYu4iGG3eU7VD9Sh2JO/9P5HxRR3NHW7hA59OTCb9sNM3ayNRW7BNWJPBua
nLPvAGD7nolIULb5zemjdGgGVtrUXhZYWeDZXCGnUfybPviapO3RyP+JwVZhBvCwyGCzh7XIDkoR
gyreYoKCANPltyhi5kIpfL1QXsRvc8eJ5h80GxL87F37u2fMfvF+Ld5aQqRrvf2pIVLHze5SR5AV
X39OEEyVKBXpAHYijQ+36Uur4wSsxnZkzug80kItgDjuxvlLy5ekZolRcWj/LVcRq84INKIhdV8c
p9raEz8DVqcA/3aHRUow7XxGA7jKuhVPut0KdLQTPAH9UrbCgRTUcJ7Fp3aLa2ouF2sNt9hxXJqg
hJ5gpQbiV1/tD4bsIVTGOdgfCMeM7knAhJSkahOqYj66n93zudV3B7taJ5iz6S75VmJShAYZVM7Y
gJyQTfVQZPTz5Ixs0aeFLyxuc0THngwHFRKDbAwkZZijSEnG0gGTdlJqIw/X+CfT+pomsIb7HlNI
aMRAz76WUJpDXWaMfdw9ohrgG/VQENmt4xD+0AnoK4WQjrb3FUqFj2ahMIe1cGzacCP07nKZuvro
aprj7WdLZDq2x2NZHoJz9j745LKorWLsIAFvI5azt4R7EE2U5sR1eZZ5/TIsPh32MMW0s64Qm3kM
Nr0x/IMyGTdkImp3FDXp6JQXWCQ8c+/mkDGPdssh4DrWo0fUj8fmAaitrPGyR95T7MfMGOAHLWlO
ivdc2okNb0qQ3BSOYsyGIkpCWXSRcsG08+kJFW0JxUo/rHKr2ZSlbCS3LMsltVYnzO9c5JB1o30A
oEL/xRABspg78oFjTvVxiOFwmnuwAwJ6YkVdkZXenL0kNBvvyssOWtOnpNK5tDYVm9N0epoD+L+9
y6ESrONH3KoxbgEwPiVHMC4SNYgOOlNzMx9fPRKSfVfxXIh0MPc4QdFR4SSh8C8AHhNJ+nTjrzb5
M9fiynoosXtB9Q4tfUUdt/cD/OCUhdSsxAMBVEicdXl/Bmt+0US1+TpA+M3b9DtAB8eY2CB+DoxY
Huu1xB0neqTyav1JoVvJbnnXgsaf+jrayLUsOaiC9LmhMOODGrwQ3m/daoDXNhOYOuK0SkVmX71x
fn64wZ0HZZuTDcjXDE5HRPSvpep7EMi4JsoFrnsqVLCBAHwHAXgv+Bz6Kr1X5Ogi3N+3aJWjQVzV
tvHrHIO8BFc9/wBm3r3w6g4dIvS0eofYk6Ovv4yqISDPcF3ZlTMjmWAO80mbdLOaEQORRFXIT31J
k+NNzXClewCNN+eWjFB3uYnF8aXWHmn5yo1AdcfghP14LW4a9LdEWUZjPUtVDTTllB7qGSbNDr5K
8INQnVFY4//oZm20WmgEPdFoe9lXi89o6DY35frE/8SKibJ7j+s5hAP7WsOtk/x3esAN1QFgBm2/
kdCBv8vXdKx7K/S+daSqIQv19Bzf5fSEvuumsIIcYQ3kGOI1jRdyA8tQpVR5QiigS7/U9O9Bn3Us
37YTmHPI5wEteFm2LI6Mn7aH+QcycW/Sz38RubUa5vuZ0QnHlXQI2Ns/A95s7FRPGbyip947oDQ9
tOKR2NM7Lo3Hd16nwETqwqtwA6luo9hj2ND8UOuErX+mTQBDsa2rtVWL6UE0FerAbCrvi+lH4RG4
lmLixQ03fk3jkDEGuoFsGMwK4GqfRqhKhzGGDJwuT+pdIf8JwiKv/YOSuZaFoqxQ2caCCjkx6M+5
TcmsDlp+VcgGKuyTXJH1zniPben+GK8MJtp1f0N2GKMIptvMhc5Oc2gYZ2l9/6jU+dV4fpEzbNEh
rd2FsJ0Kdo74TPRcEiJgbOXoSBQVGP68DrP2TfdcfPhSunrocSm3As0+Y4trFnxoD8CIq890Ue39
Gg07pRRf6O1rCDP8fdgkRdUQm1X4CJRXEi9JXlT2PhDbJH/J/oDEW+txlUWUJ597dKjjkOFJ1Bb/
+zkfbenzQDrcDkGenuH6Pi7cPB811qIMVGEXnTFcC2UGBLIMPnTgOTlxMOQimdpOviC3V8Ey4y0/
teT2XiGhBAz51shoEh1IxW7GR/QLFTgoSYDxplE40zFz5j4r4UqWhQqsK1TN/hyOqy9g63jZMupn
+w7dWS80sDC1ZbtrJogZ+t1ZuGmVHmmalfiQxc4mYgujQ0RYApdqWd7iNxOkFbm44lC8HLSN3ss8
zzNNgr9VHrnWi7KS7JnfcHL4i0gtiHh6oTjIB2LsJzK+vIEKRcQrr35XQiNjoYLTluTKtrpf03oN
4TgmuvrEXpNh6uj8H1AY+opF0e9fosx9Tu9xW4d9YxQojBWDIaeXtHn3Gx37gtbGTw0J4HddJo7N
V+aAXvA+9k0CLajVrd445z/9CditReiDDOHqOeEXa9BPjBKm/N7yb1pOiXqKmjnYCZB/MX3I33xg
zGneVhyfW6u5vvO/NMexBt1uEggGF6d2dRvDTGfkFklAe++CRPM6neQMRlTnIf8jwvXcObAlVobz
Li01Gp5x1tN3ng86ydnYjSMQ3uK5x7kY1a7NDsfK+QRm37mlyjDDy51HCaCUrQWArABryksNN/AX
S0NZtiuNrPFOTA26TXdQWX6gdh5TNL1YcRAgrq7TtJGXESuBRziGkXHZ/k7Z2nfzdm7/hJkZih3+
tla54dlLyvkGRiuEXtphJ0VDGAaY722BbrMvAJzmEQPEsGZTeE7iM19u4L4sLPckjbNOD1POqfW8
0q27gVX1arTiaqQ0x1EzKYbga/Wdnp+gOmvNf1K4syHiqN2DYxl98rBaBKNJiJUKLhaunmuEkjd7
6+UoEj1Ox515rapIGqijyY9g3728Aiw4p2y1GqCnVc3WhqwrT9j9YJm/t8W4hwQL+usbOabTuAAt
XF+bZ3ZPmfB/VFXjgcCuT+u/cZ1DUoXXxAigAYvO6zam34xQgz4svk8Jy7EdT80NQeNGRSyPcsYV
FKPsQdSHUw6gAVJjajhVGkrvDNQ8b8HGtvwzlj4qSLk6f83HKKQ18/WlgUi4Eom99TRzjExMXu0G
5be+ZBN8e2UTn1aUURvjx7abby9g4Dc7YoDg+W8MNBp+vA+4n/aDNMhiGI/JDITMrDBfkOcVT/OK
EoOouXNgcNgtZcLgzuTOkE6uTTvjBWBLV63OurPumEUHXBt29XvFGZqDkxj33VfyJH8NIGM5vqa4
Z5db5ofKRIzqQJ/ZQ9VMYecAewvReBJ8JLzD+BNrJb824XzWGwOOkshpK1iBmonH/uZIR7/SviDN
eBmU5vulfqoJFfjmDfwlq75v+ZySA8G3DuhrtcjYcBIdbuzMJRKv1QMk16wrylmO1PJWwNELN9iR
HI29E6W31oRdL8Ae1Akc30F7whB9SKSXoSWYK53kTqOs29kScHSBMu7PAoGz/fTxh/Vaum+6pxBK
giDF9/qDKaqq9eOe7oKLpIxPCwGWqpIQFWOG8SZc/48FaaaBsYSIilOzUY4RmwDX4Y1VXwAGwXK2
wrI2KhWcTL9iC3VbpW4OtJzMESNco36T3obHUxgIsX7E7Ul6F7s2SYtnGg6Wjyged/2Kaxlru3U7
5SX8cmlNK11TuvGjkcITcfyokiy5dCzrMbS2RQGUlEr+E3tgotZRvAyv3DRnZWtBLyXZpnndzyII
3VriwivJfCVHwDAH4tSj++VCYujMHClFnRri/XUAy3B8T0xseEaLdMJUtq2KnRSeGRlC3iNV1vkV
5R3kxjstB7tRk4K1/eRyy/dwrZO2mJj3iHiarSZO5XB2vz2r3ScNEegdaS68LZFRfJxjvDdGY4ZH
3cuDdO54KC0idWh98eVUmUp1kExkAJRlKGW28VqEPcOUmaEh5riK/j/LJNZWuwsZx45ssidzgN0I
SrOe6tdNVentunMVeZwwcz7aJLggoblsfpo1ba3cUYWlrocEpxNbj8yAzGSuNH5vATvNR0U+BvKx
BD2Qt3OjxNS38ck/nymCC4+xmea729i5LljMIRWjPlWM6c9f6BUMru0L7ebwGWIdBvbcuocqSkL6
KGc2AbgrW/prKw8XPI3tiicUyPP3WiksQPVEXWwSzLDJn+Ea2ggasspBnS144K8N6vnjz4HxdYDH
xRwgYHzbzOi5SbSsW/8vt9WBJ4av8/YUBfpPcx4sVWVJ8m/Mrd2lEDU/7OpjiH0MvcEaFy2/lXu3
cO+bBCeFkRvPpSv1zCZlIUj/DFSyhIh6UYmxfEBKQ4EZ39q54wPVkD8XxYLqlBEqowLi9xyCc4Lr
MNGLabd3v1gITKoOhswBlWeWHNzV4cxIznWPA/crkUTxxE8zSOYIJ7dBjzFvwyJ7j4QfVPnSiUNu
G1xPcdjH58xPFnTzbmWLVfVyb15T4sihR6HDZ7LanWxuEwsO31SEQhIJM1KZzb3ZG+0pihipsDxT
UHvurqKLRqc4G5lTIUdhPllh0CrhyDIS4yzJHr1CZSAuceZefceIQYVsw9t7Phwcw491MUT8e4hM
RiHyFDDyAVnveiMEduWn9QfIaZD6RVIA9USyyfDjAPcmC7lQh9Zq7Op3tKgj//Txevc7kKIr5KEU
y3elIGVjTaxIS/q2AIO1aM8Wh3KVE4dPVJjp+YDjqUCT9fe/yajE896ms1ATpEUfcj5uCBdv6j3d
gBrus5ep9Gd8ZLifRyU8rXSv6rjFB6jO8hdL7pXetkhBnHEnOskjtAx7aZ9guEt3BsXQp/dVL3bO
sPCINlQh+JcMNha3X8xmqHiPPXrgI8PbFrWZ7TOGmvkH2qMnZFmplXQiaqV5NXchS9tbYVuxqEx/
Pj1Hmh1R8n0QfcOoSJIsM89fmx9ma1svY7zpnq8qn/8YwlNvlBqkfDXZgAGKQ5nPqfvyR6ijQLoh
FEcjFddNtUpEW/cmGE6aYbPQZvHcOIKkUAdSj9fKAOZ6U7RdAv4jNMA2ZmELPjCxXfTVFP2rsmOV
YaoU+7R0f/y43ei270VHKI1jSl5ygyOyjbAqB6a3+UpiS7Hemp06nUFLUKPgMWhcKSd7keFbyCj3
cd65hFPmsXDaT/cdL4H0gfCBW7mcpje9N3YTVgs5wvHad7kyvMaNCU4DwaButGiKDXQkhzZLHMC5
cgO+BOPdwiW7IzKBXlL72prMfQz8fGpip+G2MuhsuK8tV/DgYvYcUkBsMWBT3VshzbIK1QhYJ2pG
az4uWxBuSgong3vQ4Xm+0e24eD9fkzC7rdIdTK71WPg3HDTMLqc0GmVuD7AWRqtAtlD1wQoKsIsH
X+d9qrote8fDIGQ10hzKfadklih/9F70j1oxvFnkRP/RPkD5Zc+wt3WpsMGpXNtkvtHD6DRiB3yT
r+5bVFHNFw0OlRbD/ZvaWFO/iaQCC4yJdBa8Wu+3+PqafsbaXub/+KvHUgYOP8VPU3oCaaKmiahe
nP/9YYeUIoROXKMB9ezn5g8KN7MPwYMOxlWGZU2zsrfOeXHCdrY8C0nQckdBDmhpHSa4mH0EkPpj
tKPWIDatecRShPuAulrC+54mos7EKe+EZis8j3vAV1GzYmHZ0csY3TSiWNnw+npt9CIMKnadI+xH
ujk0igcZYjYot2NR9n/P1OJ/rQ2q2gBEkRkgN4OfmnUowg6SBnfWGr7PKBah6ZW8j6NUPm75PAgd
mWGmKHFpkvpNY5hsMvwZ0u5EFGJy4aqYeFjCQEkmIo1t0i8KiGKO6EVNznbZ2/xC5Q5EWwLOivNm
tXgRjc+9Xl94FWOeVYSSxnJHHTgzCFpKViTWY2rR6fF6hk6eiERYb3MrAfts4Bobydtq9nxvcr3W
YAEdO8L8ANyNsZehZVSG9jWoOK4gaQOcjhUgNm50HzOYvI2M7sxazngXtQwwabh926njQSCo4+dD
ZhlYHfVusmuzrLbfpPdvz8VXZijQjIXLcxoXpVHdMLadp0cwuyR2Zql6p6q1yuWSuzqDhK0SrAuo
dZh4Fspw2ybReazgvGdZBhAqRSN3LQ8oRmuSYRAU+vmJnjPxI9TVyx40L0lhqdkF5bkApa2h09ho
WwITquM6EKnai//4xLQxulsx59EusfNu1scakGnap4xMdyt6vhqQWjByftP4+u1i0kn5mZCyE4+X
Ruwcnt3vBIZvVD+JFEIXODISe7ZLXChWR2vMEAH3dfBLRtj9vw38HSzvhg0h0mtorUmQiJGH9RUM
9g1+50YjGCpHHN+kBA6bCMbcT2+OZiDP44ZPYJjU+7uIE0xqhphtuvX4Pi6awYJ4OcFMDxYZzlEg
40I4j7XbPrxPBhCwyOhkch+3GEj+wocHG3wxcx0qhGAxacVUG4aoEiX7daLovcB00wXRz8fITMr+
D49wIeFDqqKRSMkvXXq2q1GOGvPqj9R7Uc4dyhF8mDUcMtuHD513iQqP3I/+17MEmPTFjzvlK7zj
GiwcucRae004qRdciRIrF3/RzmVlDvyBOI0Scu/U6TCqvX3Vs1xSqi+Inz4wwr3kw+Tetr6v7gPj
CgumsJ8yHycxitRwKM9FMdWskMe7XpIVBzQ6dpKHT4P9TM2tBlTWb4iDBX3E4VNbwI3nCnNT8hAE
L3D+Eh8ZXRAkOSyz7GeAMfx+0Du7Ifd9UJey6wR4VqmBFmePDT0KannwF5ZYp5z+T20Ks2JrOARV
UwX57Uh3G1ybVNw+73v9cRc1VpR5XWdEI/wRnav/ZlDE46u7zaHVngSXoH0bVM66gxZmOQTVRGlg
0CquVGvH17G1FMK3hpWCTgWL6XikhUQgY0qbAB1P1MOp8TiB/CGbhAMEx6dG3JjVjSNVTySyl7gq
Lqv9ZmxSsleiBXH81bjhDaVmc8kB20bddA0/ArxaKJUDm2pC1vXgJ0E2sqTOnNfaLbj7Xnjjynqr
/8kPVE82q503fREQlm9nuN2/sHHsHHEIcsFSxGpN1LT77MbzLyo2JhwVR/HxVJHK9RQdnV/y3oiY
/Cx1dzruG+p1f/ktFfjn0S1kxjL/xOvot2ML6l3ms4s/A/7aib4rwN6yID3e2aV1T/gVl7hGZt3W
uDnBfpoTYpMgOGDzC3DY5aWiBAN9d3jL/bjo4TZ9Rxmbt303XemurBii3Ls61vFm1CF8rNJs+J3R
zpmjJrvr79M9WgLVU6BWz/Wp94Ia11bGk11FQhsSDTugnz7ViMhPJ3zJBworgGpctaA6GIBKhPLX
k5ZnFnO5ihdzOslDGuI7/LkI3RLt52Q/mFrlhpqoOpc5o73C+RWfHJ3VGfR6Jh9SCT7LE02Qs6mT
rHhy4wBwWFhmBM44yc/KmEI127md8gQdF3B4Y8u1ys2LjaYDne2kUZKr2N3Qx+lQ1/svfgKLdtNg
4mCujVLcC+m0QzNnlR1W1SrlXLC3V3gYsj/57QKpQY1WedetBEyyYxWeXQa7ltA1c19v1OwQJOT4
E2gapUUiyG35ALknBS4970yPKXHZ++SxCGoLoO9sLGs3/ERUAbr/RMbbewMo2jGBJ3/jY7dDKn3Y
Mp1G2YTvgMSOMe735W5IABMzyhD/CkjsKK75kiSK0qDPtzPNhgN9AT6NXSU89ZO5yuWeCzSdoTOl
rYyFKVlf1iFI0EMHAvAX2wXVP9lG6W9j27v5MscNAA0XnQXirGeQjt9nsmt+2fejn0TMUDb+9v7a
3lnS4nCoEguWlJFxnUirL+Se2IhbkKxXoAUA2WLgd+dgu5nA5V++MvLzo5DiINu6XDJTsaCrQcBA
Z/NHBhyW+pXyWuYCpj97BUuspnH6ORIo8hV13/Kep5z1qIofk5+IGtmdhJdhxEuJ2v5WJh7ez4Ys
fvsAUdYwyot5RegJYfFSuPVZ+r05pU72oCEdqjSixO+ethYRptACEa0QVfVpsA0fs2lowjdlo8DU
A3fTHXxQr0PZZe3nyqIxApCyTn5Zw+GvkKoo6Qdl6Te+yylwdyqP08cLVwniuXtK+7/kWS1/2Fal
pvoY//Xv/RXXvB0rOC1eNrn5sITAYVGOaL/hLBJ30hFb+mLJqBPJmTfprO8eQ5jdzLhv+HhAhBD8
YDsidAghzUxIpX3cq/FBRLbbk4ID2sd0zbMSfMMVgb/VC2/njCjO7DTsREmRcCFnUbpwXJnso9Kn
1nABklhBHeEDuPhA62Gj/7Onbadh3tJ7dvWIIga+Y8nIvDWdPHuLVQOKITnEeVRN1tIbB7e8cLzq
c7+EfshvizLDO57t+gl6iKWfK23mhU7A3VcN3Rg3u0mtyPNx5EgUB6DTiJRmvEKoUFHwG4TGQpA8
CpJW9LqUBceZjk5hcKfKsOWFPQ/PEjz4frNg/GcWh8Zwt22Do8x2fBBJfeh1VVygHxDTr5AHDmhh
6x9AsXmPsRRbQ1Kn6hqcG3dSpd3FJe7GZvpUvfiCeSEmgTHmSt73TPlw6Ot45I4uGdrx8aAJj64+
CiWv6OH4z3j0c25mYDfzQlg1nhbv0PHBMoEH1JjrsPmAVdISPWmwbJXYwHxCLUovER/NHTstx4XW
mELLUqwlI4sXxofx4DfRMD5yuRoWrrh/Syh7bX2HQzfvoBoOcQ3SLKe3yAWyP4H9mjwdosfdH1aT
NI/+KF0Jp9Oinb+9qbS82bcsO0aT/kiAHRMrTvbyexnpr0n1s8zOANje/yejG9H/b4CrthQMXmB/
5O660TT14zoQEGo4PMORlhgS2hdCgAwo/gwyJUVsI8oARt6ZsbQmMbLYUUz/hlxcbyFhocOFhJBt
Qxp7c4RUSnw9hR216gQRzNl39GJZpf2TjrtZ40ppdbQ3wjpMZEf4yDqiitV0t0plkD1CCHrcc+Tk
i1eemXs2Ky5QU4D6E3PnHYSNllNju32QRcXUoXYYPWjhw9vXBVMII/pVrclxZrAWi0gVtFdoPyCr
aVgmAccO9BIeJecOWCiQ0euWCW/MiiK7R/jlNOrfnXGAcsMkR/w+St/7hHOGJMn+zqa9SVsAKR7s
A/kro3eY3R+UismDPI/KmrHJvcGBwvk2JlewTb1bKxnVJDex4PVLny3uixPhoAYu/ZeSx2v2Uq7F
X9eBunqH2LODLrEeAkIdHmhwRta4CHi1AAe8UK+p7Mx7uL44psFvJEaCT+eYP2mS3gJpTWx0LMor
dCaOKYJj0yNLFUX8JyN0xYEbyo9CY7qnA8xZZNlvCyu882b6vp4xPRTklbjVMwymZz8iu1S0GwfU
2KJvMDFkxf65V00s1AZNbqoLQNTyY745mzHpS7J1I1uMdlvCmqU9Ru8jIkhqSUu3oTp8BzMFB9iK
PhT/Pwp20gOuS3DvczhZscrgNmg3E4WfKzA5ucmUpCagd15lG/UdzxjsCmDIiBRrIguXiRTCunkF
A49h3XojOCafD6hGBK4UXirL3ZC9LPbuZo6TTEXNDn4vtZd0LMZSBgOoQ4ZzbzxfRVYliW/Fj7i0
DkGx3dhuD7b0Ye/H9XCOHCX+rzv6ySjM/QCytkWadmEc9uuitNULvCWCUZQHYn4uDKrQhaLsgZbL
TO2Irkbk2UPsomJ07YpH672wL9v1q4+MdOJHo0AtZcziT3XlmcTek6hsmXb9zJSgM2RNNkh9YYho
KtOwbT7/dBk1gsrb+2fwnSrvXUTc19aapfF6sY+tDvSFRsOJp8pmSwXPZfAZoF0EL3NgtxSTev/L
IBssAdPIMhPtpNyZ5xrNgLW7+ZbucCoo61Mci0LpFdqPtmLTAHdfYogj2SYlpX65Tdu8BWk8OXjG
+K80enuzesa2BoJYTYr6FpapO+YIAlhyUnFfW0XzfqOaXpIciW7ZhvZ1nLkVjczJCY4PDYoSpFgu
e9jH/HPHclqhOjYgt+UZPnCNoVfLA+rTtt6zOEgVI8nQTNOPnOUTxefE2tobBN+OlAJQBRszD1Lr
3FO/uVdCnlg1Zi0UBEIvlDoLQ1AFCIWr8GGCCcYlm13t9mVv7zNIX6gC8+C0ptB5knjYYSy5NMst
x/xUfClWfG4/LKsJ1GR275rfgUBYhmf/nezV9qBEaQT34qAkgiXCc5wEXTFx8fUZVBgmcGLbRcPi
KQte/3cO/NMNuyuSgtiZ8g25fPtBvvVkBzutZ49VFcQ3fgbDJnMtKBfnuIGiDmDYloKIBk7u9QqW
xYSESBNs3K53AoEkVW8hiatnXE5Aonqu6bIcrOqAMJK2JwpKkSlzFZQtuHimVM0amHfP4iwk7WNl
l0H7SVp0qZOne43tDKe7eKa9m38E++dTgXrLmJ4sx4/1ocVG0ZfzVk8/U4KNdExEPs+tKyQyQZs7
T9o1IRdOsZkDzNoygUHxyvhWyeRwnmzwB+wu0rRdqWn31Qyyy4J3d/OSAiIPkW7aMjVG9scBCcQs
mwFRX6/RP+uA3ALDiQy1+KUIbsYpvOFtlecWHQZzsEqyn0ZQevG1anGKwLGOs5Mnb0GsazGloX2N
OW5wxFb+DqjCWyo+Psp4Ykt9tY5EKIYoMRTCCrrpfQJ4aCTy418iIRIF6UvDUlebiswmfJuWr9FT
sWWDpQ5dPPLYzL9HpCQzuaMpP+r1p5XU02L+cnBiCZxEtflMAyyh2vHBGrG/HqaerQji6hct4Wev
lj6GTzX1KW7dZZ72t1qCcDXZXyIY8uuPmtbqQeskSEbZjxlEDy5eEagiIn0e3EXlWOD+eFBw8lQA
nPFx/Uw8TEBSLH0m/JkO1ra5r/vhOJbQ29u2z+D3ZwqONw5TSFmy4+RJsVeteNDSuqhhMiD7IJ5/
6lw1HsLb/ClGiopbe3sOuPx+gsF9sdkZMZXoUX3Cvt5U1w0LRRRhoQYnLc6bOy8vWGALSwu3ruHP
qR8We8YgFAohcvgwSrbcBEP+58VbllwOSzbrKP2O9lV7//9jcxrIU8qu7ow+hI/uUl3xY9JQ+lfE
xyIqoEUoC0TmdkrLfhgitdAkN2M9eXQ0RUvgDq8Voa07EPeKEMzU7KkTvJEQLLcLj3etEE7JwXR/
qUGqjQ0KgXt7UG7Bc54oCunCbMRV0ecbE4pkjA8M8hqwPC8pE3cmLCVEztUue+G46aicu6MWUrY/
Ge2ItByVAxUCNu07eprD3D5sX9L3zwj1BWxC4LAzb7BnFwuSQBWEIaDacvti2NXcVC9Swt8Hjb+Y
FildvZ81UbO+P3fIvK2sqHT5JIY9u5ZH9QmqPFNLteizUzhoAAnXn0zaqJ+5D4O2JqyAsgI/EyHC
NYselxYOBj3JIZ1oZnqVS1ra3mGxeMSD/elIdqBF+rUBF+K+uLgkdofd8BIsYh96lXTUf/q/w5kj
7+wpA2KLQOWaMIggwc/xZs30ezdc05LdMetacKGrf17oZxRcnH+yB3sZu7wqbDxE9HXcx2HzIN5j
u52Jwmc7/C04totqiv5m0f3Q3yVK99po3nESzi3E8biv/wLMgmkTjv2r8CHiEBuNuDhLIx+Hd03h
3tBKrdJGimusKvIZ/0eLeX3k9R6MGxRsi/55OJxa667SXhDgjz7zA0dEUxFxORucDdl+wB3EwnPR
ulsLx6mY4ynLbqV+C0+/RzvrTGrE48t6Q8oY8xBoqgyqvhJzYSIX3uEJZsUwGh19b46dOm6bHJxL
gy9DsFCW26/mT9swrtQEbbaU8kH1Q/vXSijlZnJGins2wi4qPqCjff/3AbpVA8KEryR5Yrp72VBs
ktZMKk+ag8aEgFUwkNRMzeD6416vN3pF690JNodHK12nwdby0qHZcYvLmkZdE346i3YZ+zJIcqdJ
rm5LifXXRh2puUyKYEzedmmUH37BmFdTImKLay/VybqhKcHw6e4I9QDGQckF0eZyDMsLO2Qafmbn
KIK7DjuEaI7iknpITuJMsxZ+AeNFS677tm81cwLj4/WrZI29KA2/GPcT4WHWNzQgOkCmAsfdCUsv
J1jo5CY+b0tq8FMuxEDZv3W1VgotEYJZt4Fd/hCarFKfdSR1KCALIVKeoD12a8Cqh3gbKine0P6A
vfXiIUQ+PrejX/aWD5Wov4EZaD+3nAlp0Jd/rlJSwXJw5sOTS59QtZHZ3qhHMy6dR92l36ByIC3A
oCR9wNmKuirDNDA/2IxIqzX6d96znyKliYT7tBSTVw/5PtxGwkHauNxOuwFtUJfY3UWSxHNv1JQl
cJA5P3aJyzbm9QAcwt6jcidt7O4i5kgtmjoOoLK6X2JRWIRPAzZcFetrzq2U/tfF/UgrwUKGMc/C
1mNH3XVHwJ74TrX72/L1nMguVTQJROfAvQgiIMJq7ahAgms7jQO/WQd61Zo7y5YEj+cSQMRgsDbz
bf3+79Skk0HHh994djBmnyodS4N+8BeLCnAoNolSlpX404x4Wp9+juc8f9mgJapomrXE8EvDqQ4X
XSZKmFjSnkr+5LT9Q0qaOMJ7Zb5Egq2oXEfF4ceVHFpS7YBFmbpM2yxtFBp1WjYblWITFeWQnkiv
vbaO6iTsmaUgoPT+2H7efoc6PjFVulNy4JM1KmSLVsTSMrCNYYG0ieCdIq+kg2xeamkbSpS+U3lb
pjfIYugjJYdJCavkh46hpW6DsoDHlNwZlLg9bHiz9QWqaY2ZJpDZN/9vdUHjYCt0jnQ9zx7V/aob
Pzs8AXbVmNRNY3p3jaSFk2ywZzOK7nkxczUmE634NUY81Jn9IO/8tjlyXwPFEBSrmnCEg/zLh6LN
9aEn5xrs/PbDAf3LrABSKGYDPAUFtIVVAyGUtQLXxZardxEBP4Y1VgRWAy2zVRjoXPOBPKpW1uvg
urBDoRIwPPsHVofxzz6tjvBha7wByZpZuywBxVB75ftOQNPsf9t0j3b2ESl5TGy6qnyaAE+f1Gp4
EShNx83w6wdT+kOCrKcXhp+VafgLfswtN9gZ7CWGtclo3Ah2HGwj8TtLTf5e0RodHlM8GvWror5i
ZD4Bwa6ZedY/pPWkDCW8GY3K/3YJh6FPSJ+OpGmbOZGEvC7rxOuMxbW4uU9yzU8b672EVAf90c+9
s1AfA8cYWiwXJjVhT+hU0avfKGih8WWNKr5/BYFP03u7t/hn0rk28F2gH4El6USHMCaYPARIcZ2O
8rtRr6kVcSMkTee1yKztg1EBXxuUi3h7pzPQzFIZ0avFGJRENCNmbsGu6YFvQcVMbg+YlESPgxsl
Aiz/mzkZm3X6F8dzulz7K1XxUiUuht3ROLtbRBZveLAEgvZxZcSVOM0LJrhox19CN72tfX2bvGbo
s3MHyttgr+xZH1q0D8D5BaTVS/F3BH5plv3AVr6adUX1mAYV0o7YXpuYbnxvbdE9H2ZM9tNiaP8Q
ZU5YOwv6rZPe4q6BH0JCrQG2amH6yRmwyDiLO5kpcnJ2fnN5rgItSDflJrOgKuVbXecKxesO5+4s
6gTWKFHHQdrRV3uPWuDRY7INzycSb5Aydc1PCtvFXaLVbfhfrGY9WmKbwl16uUyud5xZoauYW5Dz
gGVzEijk4MU1oUBjVFVhftZ+QLSGP3kjkRsCNInIwT4rTf4CZvdD2K80ykBVqGntmPpoMuOFHszB
2lbUeCnklWibBJWAFtlydjz9KyElbxCfV0mUuiPOAVIZAvabvkq+DA1GBOCsb+u3H2R27ZKnp2Ge
mPBHadgZT5xgIjlAOFuK14RsjXKzwBkN8vl9U2YmpCxOtwBS5YH/n8SgXxKBlmfE+cfesZUOZshh
eX1mPxtPlj8BR36nzzXDhn1Pb7aWA9vthJ/3W62f+DHAFUVF7MVLZGE+l1gm9oR+DEjCZhCj5vsZ
DIxJdMTWyEsKjrBaBsADTrbAYpUz52mrvx3XgLtVc4e7taWifP4CTgRPbRaqAYY1j4GcwsAs+3oN
7zUbJPs/bALA7yCj7UGZgJjWTN03mVv1VkYnN9mIfMy92u2SzjbSpl0xi9RJZKO9g2fIE73g/Qg3
CoW9yklZWX9RCjG3wK/kd911y4txjwabchamswBN2sMfQd8KJ5/W+Yi0pYbH7ulGYPFjXaMlciDF
e4HdpDONPjrFAT6Y3BYjLsXF3OSgQAxURkoXVoLuL6zDUBK4xgg1Zgk/SltP0LknzLwEegFaLwyE
OOu1El1MhGPZqVnq6X8M25JJCQOut52jsExjgF+DI6ThCnkDt0kYoN9c1AxOfceukq37Q8AvZLX+
g/QA9YP1nak55X5YK2XC11noZp6QWrissMycocwpIlxLkCXRQK7BDKb2THBH9BbkIVbzpVOcPz2T
jnphUV33glzQPXjNxOm7MyZirVgIm2AXTwqT9d55/njzp7k8n4x+Yhyq42J1pLofxw4X0kk5VSIa
YG9volCtUJheCxw3XKj+YwoOFVyV4dtgm0Rs7N/B6LkSAfdGqRloXouXIg4JmcNKzOxVulx25y65
NXFpZ1MyLyO6kMGP83JvA0hsKgD9JqGR4M9vosgch9paT/NZY0uKaeGqfrIt8wsrawPsBYS9GQgP
A+XjLRJFJ7kkGsGPTTejmXcEcEmkUter8BzSgemBdBgFyhpcxU8Fzw0ThHiMae7DduW4bJxuTobE
lC+28ExV3B9/FgKCD0tWRQkn5POe8CFFCZOFclWSex6WXMzqp1Lzptqb6K/KVyQH+9KYHfnf6/iO
g+2V3f76C0nfd3ZJve5Hk7bcOLI1pQmFwqGSKB/OS2t4MWtEFq1sLTonNTmeknhcAP2CgX3Yv4xb
VokwdZjvZRO/9Y45mDsUNogFY1g+03+TTTkwsd3pIkxWjcehESCroSXyEx+iUtOyU6qu56Dyh2Je
UBCBI7OscFQFSsIrHJObLKXhHSwNAJZzU1UVQfInynskFkleV7qQFzQhQ0V6PM7BnUuJtEST70u/
VqcHCn7fTRH6GFVPUqUJW4O0MW58jxk91T5JqNK2pigAkd3o7R4IUHX2q5VRCmgd3sDkFSdUVZUC
tWalpy5iInXhbKDeOXcMZJJ/MmpeAefky36Mk+Z183vbyspn85fOz5LMkBMULOJgFc4/mPJFaOgP
GZhwBNXrKOMkyjOwodkBFLmn3WAMFkbZFzsRKww9WxwBqU8V7goup84CRZNkij+LCvu0aQ8vu84y
dDgFb9oFQvPPI5MsJbN5TYas9SU8foOEAefRQNOGT1/7NoYqCWmT9bnpf/ytIHIV4betnTc/RNfq
iB7XET/UPfAXRMXFZTq/XkKFbmgmWr9U5o62yTD7bvuUoPadcEggcHhdPnuxMhaq6z2e7yHQbAJN
vy8v7FG+X+d15dojmPvzV8NZzcfFhVAa54c+7XAncx3cm5mkKibMpIMXTUfMCEkJyqujln/3Hslt
zSFJ/kPnEb9uSurLRYjDrrQMd+7bJvlLWNSGm8BoUN/y+K9P/I3SjnxLUUm0Jqq2TQGJmuXXX6g3
qA591S563oFEdcRZ/JclnLScgtOQprPYlfBpoD/Sfo8OzBPrQvPSMQavvlDxdZxusUAcCDFVXl8g
NdqpP0BzhgUr1Z3nY5wVsmHtmFxX0ZjXUIYJZeSaas5nGHHNTvVx8/Xq2QyrYKge5g83sc4oOq2+
DmgAIQh8/o0alg6IBWeYDIZ/hS8Wb2+Q+eLQQLvgF5esFnycNmd+DUQx9PIiLzT2kOArK5+WV66H
07wRSDxM8UU5W+oEFdJFFabt6toWvjiQrpij00EjOI84A/ht6mWNBBJyaU1pTZ97GyWAVCfg9pLo
lzTxrbgsf0ibIkiozZK3ZkR9C1VjEawoB8NKtkM5QgN37Vas+Ua0TS2E1GddtZ3oZh31A5hN8DSD
KpMP5dFER+YUjVlQKeY8oMzNBnClHdi88Er+S6mkF0pYRdcwj64DFmk1LLDLBcRYDZG90RUJ0q7i
Fh1LkNqITW+XEUdzTUecbsd0gZCJMfj+atPUvJWQ/u+78WMDEqUDR+JhwLhImcXadQ70A87l3zrm
9K+xQzcWMsPRgK3mWeCcD0VsGbz7o+CTOOck54cCTVZaUS6fJXKDbBJBO57ow3Isx8cLSrtznwKw
w2NZTMNuagc9KmhXbgAgB0NHmDaJfpoSl5JSvzzRpapc3gSnLsIYoHf2m0VSzQ4hRs15+uGI7gM2
e2e4Umq3PG0DUxaBrUi00vIsYJsETk9SMGtkhQGGjXoysPYo4+zTv7rjeiLfJtm/MARKhNJ9Dq4F
3sNMTqsoS21FS4NHPP3F3N46YmkMc34IsES4g5e/kpZ78fDAcWxTDp17VDrLlU17MepgEDcqu/B2
jN0SfWJfVzL6Jqk4dBt7DWJ0AAvIWFM2Mxjx1Qnui7TPdl7qwURwO+B3dguz71rDr1JqW866Gfnr
oVbZjCpVKHa3bdCW6ARoIP4cZD3/n8EGy8s1GiI+cNg8QG1C+W40zdh0Vw79uWOzf6FDn1QHRrl+
FSR87qpfjPH1ghz7EbvURU0va+8DoOItSwbhIEf+f4eVs4TEIjpVfjzuGxpYli6YiY87Pl0To02f
AnVGx5VQXGxk4+z1Otd3xa4Zamx1Kg2T8B6pb49r7lwQi4SanB543ZOGL/X49fw1MTWFdZfPyRC3
ogA4zu82FD9muVigRuyqnQ1I3LEFlXxq/nWrB0bRlkwSTqcf6RrPukSsCt0dbp4z1LXhgyZDJEfk
X0xQgGe828tF/eZGu17Ya1Al0JjyIH+qVRHOl6WiixtB+aNFA/Ar1pY3ZoG5NySLO0VMMnAunuWu
zJQku/fB3B5D+W8iYMieVMZFe+BKA2nQpzIuArfI0duXEWBPf6SV/8RBkMFCXViU9OuwWjsmBVmg
Gq9kGzxEZVaSSCJzWVl1klfLweBf7t0gjRSVNmnfLXQDjKKJKJODaqDiQgaMLOxgCOC5VYLSs8ZX
k/Zd7nvm08IzM096UOdcCNytw+SdE+sjwGU2hiu2LThdW9PUJGIMUe8mkMwAzsvXlRNo6fRcYVt2
5NaU+s3Sa4zUVRo1MzGck4pb7sC9lQWqwKew3YZIUgX7OWxrZzS6ZAvybUn44gLi1IQTxNCSun9W
Yf3Vq7G29/oedr5zscxbUM2S/t0OGcr6/xLnyDfJ8XYMOxTjmj3syOlszkqHirgXA5DUQk+4y4ea
vLakjg4lM82MWsyRp5aOz5pwSp5qO1Vh552uFRP+lRU2RH2RigE+5SweKbVD+2hg3b60yszDTU9P
xoFDkdnjHuIvOKKaguxgXnp7GSScOcdJyRywPciVyB9dcKUMa+8A2VvqFZ8etg46f8d77GQVBZKJ
fhnKthufJKRtxxbvEw8Jp27IiCT8ttfeGc4zrnjtlkk8Bmja3g9c3ibtlnjIXHBfqfMVLufCABUA
UkYqW58njufSaVMkmkaHFBvcfNW1lytZJojhBAj3tnODoW2ou1Ekl3mFEsXSb8SMmO8VzdOMSTwi
h2Z1kLZ/eBTjENN4B97fqFubclviniWIp+9AaCoqeahgqicoyt1Lt/wtkFh6OMeQCSZsTbNyW/HS
RNFobEmE7TcM9Z7zFPqGnHuH1lbjYcL8jy4TYkTqfKjC7C0vQars5qR6Tw62j1lui8g5CDp3ONNU
E3rAL4AtQhgTaCyFDjtMe+lDUFV4arUOS4QDeYVYIu/yXlkDzWr+lckNIL0hpcnt9U8QGOKfGpus
pUGSqyfG8I1rflpOcCzlx0agRCV43nCbwLk9LpG0H62W84MmrjF6G09BJKiy9PBKPj6TmoDffCZh
uGACoOVrSaAG75qI0WhUjiIgpI/wu9S/CTLb/jqep+6JXxWIjvqyw784ecBqNH9gjogA+7jehUic
akJPrbOrPzZpLj4yy8/7Vr1y/AS1uzEUsFEe8NyN6nSaoBxB5xWSqpGRbG40IueJb7z7zKKPbq1W
we5n17EzKwvEiASag4wpbVuqfyUO5ItmnmMbWIw9sRv4dYZfcH9yfE69ozlocif5UKLUXAyIcsX/
uRSSkuDJWBTP3qSJ4l/EavXT8+q2uQEARqqLIPGoyQVH8uc1CvhMApWAra4zzv8dM+WDPmqetkOB
my4nHInqAhHhaDnQyAiwbJa1NJ11k0HtFTRMHy/MJpBfqrefP5DsmqGRclORh5vghDmGPTmH2I9f
zvakr4MfOjRzRcSpd+jBC66fdp/MXelFDxTsGINg6Nf94Uuzwq17M2OJ7DNJPUn/Qof7/tRtOSOJ
kzeqaQa26RC07hjyYz1iqmLj1jQPz/23WJbNECZlBVa8lOIM3z62JFVmfsEC/vAtgU+2MJ+tvCMG
95YaGGxdXn9aRrtwSmqGbJ96WFGTPaRad9mUfC+mgEOa8Fy7/dlNSM5Y8j+HndwiAeubmg3bt8al
N84xvAufGG4EJ7TGsaqY4M+iIlEJLUnJOvahijjM5Wuv7fvePRzFkQpWgFq4XJ1MWqrFT2ER5TFh
cC1a98KkmxxPLfbFpm81e7VqQsgkAJ/SONhZTt9KOapPHp/xOX/DwTDY+2VliFaKLHbrbCko4bSn
kqEa/QDpI77rL2kFEokPOD2eC22FwcZhtRglF1lwhFayfvbMNo/UAHE5Ae0gKA46WMocoZW7sJ+X
py2Vvxt0wbdXltfP92ZQACvP9Kz/gke8ksVf03CVjsR2XPff6tMLFunGezAeMgxcERl5G8/wGGm2
5P3e4EBZieIzXw/DVJH0MIWgAuP60rJBjkQ3baHEHMW8k28NvdvpDYAGjOk7OgEKX5ZwpbCPUxhx
DhV7ZjxJa+DyRk0oHSvnwKfyf4I6wH2F3lCTy88/JB92+EHSOp0p0X+yTT+b1Yvwd0RjFRhMBW2j
T+BE6rDuaZBpBCnPJyWqxivAkmZ3v2r1gWeyro/ANULwzx1Ixwrk5ikpTPjdX+AqMNdoXdgP05oe
Cky/DdInrsUDTjMpRNNYiG8unkVSdMJ2bHwb6ySjcghL5cTBJ1KqddnTngynT8Tmon2ueN2vln7e
OGJS/WJcMatL6Zmh3aO6MUzrGIsqu4mhiaMcjX7kVe53RsSOl5Pgwb1Z2hDTlxgJ2wlmD3KA3vDS
YW1e7FJmtaeajpsB+OzQXYrpBrhWYfC/+tRYyxewOHnd2sz1QLLwI3d+g4MhYuhe36oY2r7UQdMT
bO4g3CiLV3CYKXV8hyVlIkw3rQSv0OnW5x0QhOkf1auhV5mTVeZH9YoiYrXvOO9efKZ2GS7b/QeN
VEjmO2HiH5R/NuM/gVrmGARy6fleGEQyr1YQdW8zikjeOdp4gEJczxXHGh6fbbb64jJpkMVtG9Qe
OkFEV26ZBja5H3iHMhPnrGCF0LdhzfpehlACL00cgqPIb/V899Mjg+SlHCBfE7jZDDKPSRajHx+g
3WDnSyP5WX29Lweaq52r8YnENh5KkDW/58zFoV9iv4B95nxH76WpCzkaDRaFYZMl3UrYqOK2ZS+5
/4nBLoG1VOU71GEEeds/+vXennKawPkGd9QIOasI6V/WaZPmyzwFK3EZfY7tEaHsxo0tndnw+YWS
6reM5ugr6rJHTD+hOvW0N/bpseTuU/lDGNl1S7okLRBEtyhSTU1vMYsFlfoTz+B0wlbFNh32Xl5g
LoIlrnpSnFjd5p1hPPzBdc+KBuDinpoGNv4KAkLs3CnAprGQfgn3LTaUMwpOkTIXBQ+QH2KNmkWU
b1FYWlN3pwpu9VQ5QLPTP6CoSXiuXXm2C0aVAL4SyoawO4mR7ZAsPrKBm5c7Gpnxct/54+skleyc
T5LpSJmyP2bQopmelz9jLvl6bglK0fQWuSiFO8IoVyfoKi0scPeHne+VHvJkRLdLpEj+yP/aHXt0
kexWJYbj6Vv3ndtsXpkNh8gCHMhvFM+39tIuv6PA4K5rB5S1hpKlzXYYtwDG0xokQRf0RMdAEeY1
D7St/UOJ068zcdoKpwOHqpd0/TXsecvIWJ+vv5CdCMC8eYJBHizlfuJFhkPykXYkKdJWHWe+po6F
jN1fGHaxuPegaGrQ1F01H/4OXC+F3RPl2nX2JbU18NTqjKF0xYbjvBBoJNv37UBZnMFHi4KP2KQF
r6pzPJm9xg9sxsI/TEwcwQVeAG86WxDI9EoN/lx4/6P6/kcUVU4oBasuW2TYwnh7NDzsOvMi+FQW
xfFKJQCzFhRGmYYampFsINqaOqt/prt0BPEvqk4L26LU5+M6ST0cVliQT6F4KxM5Vy1CXY/biM8I
righldC511rZflHeX6U9lcj14t2zsjwE1JS94GpcScxM1gyXwwtdb9N5Mx3oL6dMnSB2ih8XQciA
KVnrJiKcXlR5X0Av3PifIPdamAYnyzpmZ9GQ8fkV2Gwh3wz93qcSl/W3uNbj2nXB+wu2KXxG5aYj
mqxwBnZcnqk24TUtClk9YaTKwE3/fDHGNjs3z64QljiJ0ypBGvKuuy8zTHlXkhF5m167O/F+utc2
XR4tr5jv6RoXQTI5Wu8eP4mDKTFfA3pRsOn+ovs2NJqECpwr3rvBh8iCmLafKFZNgu64FYJ00riF
SBeoAds9gmLcFk/a+hCfExqP6G31HyDcijtnPIkb5CPXP9r7xaPTyyQD/GfOQPktf9SLptl+fRUJ
40mqR+H89HHrcfLGutQ0CsA7swpxUAko3G8PnJFJHspvj8RAY4de+EQ3gX4DmSZBYAF6TpCpdHxm
thRPSAYaUcDufx371ZOwt1N7zibTUBhPSMygoekgW6VMxjajarnvvBOE305gFuFr+eAfuRw9ANj4
Wupu/AW+mbGAxY5XWwcTTpw25NjLqP0dJst0uBHsY2h5K8/xMbobncjJSMdBIrdbTlONj5MJgoBf
z11Rbmg+eMVKmsKksCI7pgTqTFq8s5PyKsndWWgOsdSy0KLV3T5jffdT0p2tRlcSIU+K7XnPJ6J9
suBGMkL/te9cRV7M2rNNwc2hpyspirahlcJhJnExA1zhi8xQNIegq4X4dhczgNkd8dwt+VPrqEic
iNFPeyd7b5R2OhCI86X/AenPGYP4eMDNcBHzw3WEmRyDvs0BayoqSZaimYi133E2/JEN+ESnUSqB
KkrzeGzJWKHcGpDjF58aAYCf2qllhScgQr0Jd76if4WyuDmdMD3QwZKTqeZjl/ei16Dni1soDcFv
fpeNEtAy8AIoyhosikdB7Yo1mXJk04PN7VCxHct4r65svHIG9qbcwa8+3QBZ7GK3ikdohUM/+34L
4q+M7FjRuuFfcV5rbOz9Yvc2I2IarI2dSMlDR6Xdu1/StptW0soeKo2nJzYEM0VPY45kIqRKxbzn
8kFGf7+nbRQg0Tdfh8PxaRYQxNDjn/JhSzocj4hCS3MFrNDErsA7/FVtrZNSQY8B2t4FS7BQ0lLG
bWsoRuixON6wKAwriJj1ktWJu73ioU+vUiJfOe/m+ltQHPOejWjIXnKtUKfmcsOPAk6syHzUJjWV
nCM4uJnmpU9T1/yh1SKBZ+rb/uoXqFhv5CHOfCSpz+zZX5QRK7Jwt5RV873W6+BSZLk/hcXohnuU
bP20VHwWrjLvi3IPGRoVrSeot96A8C8TbgXbrGPP5rmtrXbhLN+XxZ0WcE9dNb5xePeTMbKMEfRT
AeRFo4lW/Afw4ZVKA2ljA+kPOES6vTa0HiM4oPY4v31JEbbRf1z5Hs2t0qWYtGwGVUFLKF3b9ZX5
UEJDxfXB9zXBFxQiQVcTlpi2s6Xo0QbrgCUCb7AJzFEO7Nk5cVus/5pZG1X6uUTRTFJW/oGAkYND
5C/29r/O2/4UqHnui0LiXaGv4+vvAq6CnpnHldppYtSxJS9za2f88PXvbtcgDQAlYt2vw6ho+DG4
Uq7O3N5NepN/EZUmUv5J+Arrv42D30+pJZNsra5lL1WcEJI3rC/pFXFdo1jNz0INQ14S1V1KNzJM
iyi1oYWtPsn4ECe2y9eN7KCZhDDyk6+Fb/oOosFfhQG7p+EmFt50Y0zc8h++q5JCqiUwixl1l10R
DBSHpf4oQqIGYpzBqfWjxxmd6eFAWeEhxUJZFvp7m5UgAjB0Kc4wgxvS/dVZOkbriIvygpQr1hjh
mUCqbjwVw4yrhzgzznQOst7XzFHno0y5K3YUPhO7jL1KjDly04a+vtNr80VBiCZlq2ZcERZX0CLm
jIgHZTfIKx7Hx0LvXqODCCOmlnIiW9WSuvI50PIXVCB2Tcgam1dR+2Te+itSmHO7pSIqK444vpZU
fWkn8yEZjyNzh3NMgXawAtfoui+xQOYRicMBWHT+Y/6pTG1+FyR0IpUhYR168iTyxvsuHvU87ClY
m6vdJGLh4zuxtgqvfplBEYW1THR3ECIt+ISE2fc25rw+hRH7C/Md2yDVmvsUg6/Wca6knzn1fbDG
d7Cc1qqeRj8w50pfC8H6ssryXNMqDzF8YBCfi41d6gyhcmhVlYeDofSNXbH5ltzz8upIXbKh63eR
QryHKC3QgrkSnqH7TdGGfEHSsKiuvK5XND/N4BgXlBecnwNBph9sNIcDjHievvn0H2W3Imn3Ghj1
PJGHql82j/S7CvdVxAo2jMsQKtFCF/0HbjdPlsud43g/9/XK9HxxkKydhYiIK8G6tSgzwy21vbtv
Pyho0vadejjAKo1MNJ2o9zL5q0sr7d4FczSN46XlrCTdJ/LTyPOQGtTyRoBmHUiVIqy0MJ3c+mto
uvzt4Z6M7szkLPAF1ziP0Z5eA9mfeMGYDtqbGAc27sEOIXIiY3bvrHZkykefwvn6cpVFhV2wJSDW
zyyEN0ZfzxO+dZbMe7eLbyLMhddL1Z31CToRDYuGdraYIc80TVgBqLzxPtOXAlfMM2geLGpZskHL
VS/mduhuLCZYq78zeokqBFCbZ/t7gVrKe7YpArCS2lVS4FIY9bRA1+Vr74+a9wUT2H/c+8G0q6Y3
2WsiWIhVvz9uKRdQ8jJ49RfZ1HK06UxVxJA/thvycfjILJXG5mDQM9wldOJWYM3zPLSPuoJUgDH6
juy3HiGCUEUVrRtm+wRnE1lK7t3V1UN5U5mO1vfwtgjqRfz0sS/ZyMnfYpKRe7JF2TBUOe9lKO7+
Qlt3SH7+qfnvgDNQMguv2R45G9jzQYunH168t9C4/DclMKMgFDfl7S8j224BKh45D9FBbuPxeOSS
XsqZn8DTH8bq0Kp7G5jA9HaRjxF1EnoPlASWIbCg0R4ZRmqyp0eYb4cX0bm8A56sjfMDFswf/+s1
hrUqY0Jo+LfXnyuflJqiV1SWrC2qf+BIwvUiJat+K0seeUKiLntc5a2Pp4bi9WzL+JHOkudOHrL4
Q+tNdSPZbsl0WaAIJ+AdvVDfCuDadlPvqiz1eiwxl7SvQrtcyHzbZCzpRBtDM0/KXT3z994x+c/a
UpDph3LP3LX0V3CwHV8soy1ikRAvN/iXKNbUym0IFGQ+4kloPEfPcxQi0N1Ud+aGr+eqmmA/+ija
9PR77NYEpTP3suSFROQppXcpmUexhkuI7L5uGq0y1u2O+DFw9/mc6zaD10cyDNeHcadyAe8TNfRg
1DucysqAHjnP2nrRSumae0pS50XU3+Y8g0jBvTEhFr/5ObC4s5MuL7ck8cTzjvh2KD/6lGibYPa7
xSXP9YL+bM/kvZJruLh44B8nWviOep9mfTTUwpNVsyz+WEoRh36Rz8PSSIVbJEkU81TLb/wCNC1R
mp4i0sLkGeMcWFmKq5uplVDeNMOp+mccVjXqBjIlaNscaw7J3i4VDc5rfv7UHY6YgvuQZElahgkw
1t9MOtUINPuwv8IlaBlqlQjGhp0gCCfFCoZMydbLtWM8q2FYp2vY7wq1Uty6zNbf8vf7QxaSN1Bx
MgCjhb9qcV4HKgxBZvwQzLtYkFvDDCGIpb/g+ed5FcIyd5KGOY5aobhWlVQgiun5C1myInX1WRR4
liZE+7Tlizc5ZYH0aPi2jJz9RNuyInQYcyUMux6c8bWzn6XogOV8WjScUrIxdls6vkt5TZlgP7+q
GmRQCK8xQWjHId89WHXLEpfhwzxXFcSgwcvuoB19Hb8kqGmFY8RvxYAt9iwhr6fWd9tOpoqTJvtA
rj3SEEfBpN6QPsnQ28/5QWpdQ5ShLAskNrFRq047X4CxyZdQBtOzOXwTJxpLEjAS1IiLLzQEXpCA
0F+huZi/fmMsdSnyYzgiHi1vTjYbjUKelEnxDMZkYpZKIABJF58RLlVmuKzU6ugiKRu4cyBN1Opx
Y6FlYkvI/K3Z4lMHXoYS988ewiUsxO155k6NdIdi8G3/Yk1xt5rihT96Rw+w5wbFa2WNMIO3N+bm
L4ckbdbQ3mD+NRo40iCsYYLgh15vAEV0vz6DpyjOX8xuo+CiEg4cJDKYu82e4QtbfMd3Nj5sc0vi
uSPXmGQCXpR/+Gf3VG+7wLXJXCBxgW8zNhLpM1ONbLltQmzYqkuYggzIOF7AxCgEbxSMTxu1BS+p
+FH1NmRkmyBJNUB6wwTYbWevZaBOCfgtpEKdgQV59xiUwCUS5H5IO259K6fHXWzi7tudlvpm246K
b+cPjQ+bbN2lfoJ6Nt75bmmzrnUATbkbbRtsTwjhtVEufECYVVGUc69Vy06ThnCpQquAIbqr10nk
C2p98MuqV3wpIDhpQVHcUrfw1TqHm7PZNolOlNR58bVWR9d/DPEWOXLcsMop6UrYfn3VdYxF/891
ERySO4b1NSof6wugtjCn/qiBAzb8x9GA2stYlhmA0c5M5Oh4ZhqS5A7HuVDIUDpAFklm/rjtvtzO
L/18VSx1PgDCXxsn5lOof3Ami2E2DbSj671zoL7Re2NAvwWOVXE+9Pi0E1R2RbsdHKfeEIV5S1tS
A7JaYVgaS5tdyCcto1xEc1UPbCXdey09rzAWYIqvzZ69ll3aVcUe6p2U33mZrbpT2t41lAPoTyxc
Jv/7uJkXV0JslNfuYiyTUZ/8v9/FZhZfMsFMfIQGBUzzlwUiAhdRNYTdRTURhq/4qTP8tYwP2w3p
gbpXA2ZIFfSgo5gPqAgNxJ+trqUI7nGGRJaiZEHxsbCQBRkXF2HnJd253UaeH/yx7VuwXgOD2s3R
JZOf+EzqLhFfUm1OsmtDo8V3gI3l1ItzTr7J16rllgVmB0xVDzyRzs9VcuoPYf5fzR9lLeiBqLA3
PHIhwvtLomqSQhueVZw57VrOpfEKgiO4NN/e8g1FLGcDpXM68RI16hpn14lrTVfvJn4ZcEhdxcjo
A0RJYxn67ljbF0P6CYJ2jaN4w4tIwLqrgD2sDrDIyTNH31wzEnk+ZQjobNk9DV7zZGqYy0yR6gIa
qZKY59cb7VjI37uOM+JPMXIydW7CPNfkVmPyB/jZyLkI8dbVO2mP6woVQkC6TuwPqhSiB5/zvvOG
sx8SxMD8hL/ytB4xav+HK3QQJpk8uklvRdiiQTENw2hD9c9YtPniEHAFUU7Vd/LaySiBWXAZOoQG
sGAwHtxA9XFf5vkxlmcMGtfw0zGDZ39WUTFU7hM4uMqoqS/2rruutyfBW8LiSOE1px6tHwH+p/Nd
cs58f5a7VWizlqcvTpM8fNU6wPPEAgzEXhoM10YrnXj1Dyc28gmxka5FKzc+z+w3RqD5SnmiJ1y7
26cNuTgX7ueEMUlN5rCG0hM6vXPH6Wd2CyOb5JfUWNNyV4ixBswSD6FBOULTqwZTLXS/uZLn5rDM
2LqDYkppD7vlg5hvOBqywgnGJtuvCOB78+YYlhhHcES9quz4sfWBUFH4ZRSr8Y0VyHJdXIEha/EB
AsPB3f1zFZmKls0oLIGvAvqEL2sJhB7oJ/Q1bkwdBiG7jd0fs3aOKPWoh+t2fFsJgskKOZvCM8se
v9Ld0DRDwoxQOOYwKOSSOXx4SdqKESrQLzIgnvc+ITc1xxhq9tH/K0o1E5biUXfyNJFEzKxo+fbh
7dH5g0/TYME2T3yj8em2gbsL5d0IgYlRQEY6sgxOQ00nJ5eMF4fXmsvDMVk0H6ZrM6gwpOsKJ4g/
SqvUbeAwEQS9NGHZmLeQQXl9jYPZzh+hst5iPBCSPJkx+HhgF4O1D7oQXu7fnTXtRfJYdVTZLlEI
cCnlLXpx1/yfqs6wJgFiXnmkkUV10obWobWAYEQrieaY/6arJwDcQu9PqVVU/rr83EPNsntSEYfX
DfkwldaBiseL2XwEemH9cAUjKvuoNxtunqpbONpav5n9jy90ptQ6FBqeEPPWAtQUCfJWU/7EQ7en
NZubWVI4zof3ZzavfR/ROz5PQZPN3ItyufuSFfI9QCLZKXBN8Ohp1k4CsFAzHGcvpKdxdYaDIgRC
nTiNmKpvnQVxd20v4+6Cvxtc6jt0S9jQLQApoiA1Enp0EygmzO4b1yQRR7ms87NyGX4FjOeL9mko
47XWjZp81OtBJ24mZjgRiPqEYi4KDEvrJ6leAM0y2BD8fJWqsDFbRugvo+M1AID4RyupWqEm9ZV4
CB9asPgDVWERTFZTj2jZWKduST3IASi9pP8CLq2y19Q3xefkhQkVCF8yOaoz4J0bC5HRAMw6HRHH
++iTMalGiWN8+ETMf4HPpp2vYq6nZVMiCYeaiiXP2K9EzHAuYD+VfTTZxirFjCvJeFVDWPQSIyfY
zAej5yTaxdrMrcdFQDeOG+gmqRlxCtlU2RHrDa1xkWJYIwVvUf90fjyp26ocfVi74RfpcId7yDLL
8cfSmVYKwopPvDqVMOodeMM44j4DtFexr/e5cOlui+KyjAQh7a8Tcrz9+aIXaWpggeDpIMDrCzx3
Woet/qxj+NFjvyiiJP5OrqRcqx0GMpxyXDSHSvkVJPwJOc9t8sPuvScGz0Q2TwqZnzRq1/A2R84t
F+W9pCsfP6qC0rHzgyx+Io6Mr0qcaJ4TeaZkBjd3ckgUiguQoZpw+SseU+fOc1Hma/nkcNhXrwzI
q9R1ReIUTx9TI+BqDXLstyznSf6sGfbaINBJwuYpAFkeXA2+c84IBnGyL0MZUqf+uDV7CCeR6Q6R
rBdjJlVYgD4temPGbIMopoL4JdxCeNpKtLGWolFJh+sW0d0NFoyU8oyR8RTkhpbqY4GCONhEptzZ
Npd4HR83MzmvUsdYSWmzddOi6ieh4a0kZC0iBzswn1bpfnrWk3OfZQ9bYuiYOlFQDnTTJaXlEZDm
qZNEv4AjLWSyXsjtrmHsERxODaOj0WS/w9kTADWzyfPmbfxt+OVnI6dn4BQMMGsVIR9hgxhc9s48
FXPLMUNiz5z/cEn1PACMOMH5EjQNNwD1N5OLsqzyuKrb0YBoTfiU0jNE4pqkmQMrssebs59bHycq
+wHkAao6HZiBQUWolxGlslEkK093lhfnbF8DWGDWHVfFZZ8sRjbCnB5AXAtb6wKqMdeq/csRwf5r
q12b5OVtOl0oNw7XuYv8Axx1KaqBt5vQ3yXzdxSafDK5x16WxGn6pajG+I43an5o3+UvXJlJEsTt
r9SuS7hPuHcnK1sKEStVMojw6hjaTT1XJredzBXQnqXVYGUah3hyUzD7ZdH1gU5iSorOtAlS36Ne
i32PFSwibDVo+y9Fhzoi1BFYs8ZzCeZVALeXwMUMVfMTZjB3Uov81Rsihr7e4p2FjeRMZlC7tRe+
h1+MHhXGLlnZL5I9X9R8GaYg+XOj1bw4rHzFEGKfqKiLSTWKxvF4ON4jVpEpaPwEiGsYvwT8QvWY
PzBvs2k/9sLS27+bDcFWVIKG9b9sUFiHTMZiqfakVQMVg7HXGwt7h1s+l50dx23gPKW0S9FIpKZ0
Ao+RJKF5kpJ2qOlOqWmaHCLfIsw60f6kcBW4DE/odP7m3Sjc2U2TVoKCG+7k2VMHK7iSBn2yr+py
BrAxsYz6HgsgIhf3ErNz4F1fx0qV+4bhkhf7+CguSQ8X1zmf8wJj2Pgj0uozskFsUa8gWGCzeUQn
bhJHRCOjlCVl3KeeMMCFAAfJsmq6cmd4mRiYUSFJcA9rzLO/VbVpUWi/D4akPkv25iB7D9VHEo/W
fUTe94VEIhX/xZQYitOB5/0Oa1FfdAKkMCFFN6MpG/WB9PMPpdDHWRPj/hKbcZzIQCPuwuvwvNda
rB2574CH5xSqUax3zTfOJKf23dt3kJ6F4Un0aL855w5LrpqecWav48dWO7eWflZj2FSifq8LoBhy
bp5ucWKrjhj3gNdMRHR3wEyBXNJFfzEcbXAFZLSDiVRbBSDvnTX9yMHhfZrPZ4POBLLjxIXWsyGQ
bKU0eiL5tbTaF/d6lXV6qQxyYnY1eKoDFtLA7miLQCUBIUiHZHM5H7tQA/6yATj8n7u2VIIf7qeA
qOTVQqnrNy8eXcX0cP9iOAaTPZlmfCYnRTvmffJ/P1T010JUdLyarzszixvdU1ZhiQWlwNDz5yy/
XKmErXMyOa+2mAZ4ljg/cGEDN1i2iwABB0JDesc8xxOt0IfsAP8XYr6myuj9DVwh0wy1GL7T1xKd
EMXVPt2hg5mmxTviScBYdQRbQ8i+fhRpN/TJ8joI1hu4GOb+6rroU5c/anBDhkxGiSzQURpAekCq
kORHciqsCmH4A/q9RPmlsIc4Yzfp4YUrrSIwj7KCk56T7dqA67rlvvVnFTFlHGkcumzInTyqb0lH
7udZnQnpqdcBbdIL2/KDOsgEFZUM1SZXAgSoSnwrom2vefpq2pa98yLiV+bV+eR3DlEY3skW7REO
rOVzBuJjb0RUeac43IrmRhxVwJ31orVFZYt1a2DtnnhvjntqKvLXkU15vq3wrnt02AWa/nAs856h
HVaJS9zrTwkEwC51ygmiMPqVa15tM+UM5YX14xMz+uRC1j3wEQBvCHmjK9UUVdRjlOAdDBaDQi+o
t5+P8Tre9R4rbX4SpipvqI1XaTVouVWq1+4xMIh0qQIQ6l/SNM0MGu++pUYel5Y5dXZoGHIK03uF
xB2WhyG5YmQlWHym2jVXJO7nKPoLDy0FQ7SZ6ovOcpmDdmai3x6GaxZxPGPlCqZLYRZxSlcQJONH
mtrlt+l85B9FpTyRs3KDP8T+eeY13DoHXhzO9rRJ4FI6jYJYb1RzrviGjd5gUk+zsyalv6qX1c52
T1Be8E3tXgsvA5r/uJN4mWzhL/aGbNjJPumkXSQTMhuE9jFkkxs1mZuW51qKncWxzOwNdV0ohSOz
FgefAHzOTByCVz29ILvakR1FzVzTTzhepoel3t/6VjPUb8ZN3P1WrfoJt/tg+Cpj9WF+1qmLol1/
NKlaUz/YS0QNWXgrMmHpj3piokXbuaGRy5Q4VomJWdrt8yJk7Dm7/PkMixx9xf0+TuYbQDAmN1uj
aouy4sf9PJm2U8HGXV/9uXJ8sU2nNJvSbmaK0zyRtg/1YOPM+xWV2HQzR3uI2KcS73w0tSBm/PgL
g3tPfPzxg/1kXGey6kRpd7hcQGU+A7hDaEwfrgIKKeIL041PVVvmqQG+LO5sEHWiBBiO8Bxs0Fcj
Xxw9XHCJqW+mimcdrKqJRGL4ILV9RaydGNC+rQD75BR9tY82NHQvajT8f6ijpnmV9tN5T3l2SccF
DSH6C6qbHPHa8Blqn2LbV/m3BRunK54Y8mYj1BqUDZJ2oP34ieFuh+MlDgPuzasNSA86X/Ut+vNE
oYoFIpT9He7J5uVniRrBT6spSMmIjC0yhJSY1OwdNuQ3J17iolUg9QvbW5NaLjMzLz5G1Qp6DMST
snynW/WRKqBypb8b3O66slZoAZ/UzYqlK4regtCpm0mTEi2EfTmlcPoU86b9fx4wd7pFS2sKehLC
6m6zgE2kgcMyFdYzICLHK9toaEaFbKF9h00i8YRW1k27tJM2pcCJJRlp0gZhiFfeHmrL5mnBv+2O
0MBCXTQdW6lu8rpPhoNeTsFURi+8gOFYF54yLV+IaLAUZ+zSQsM0GROF7DWdb9vXloja8Ky5tR1U
wc3qjcDYP7c8Ymv89PhVBz12kbsafRW/c/jyzq3BybulcRfHgmnF41LhcD1jHgNSWqFYYrvELNEg
4XgdlzGPC8rlQhcV56yGEFdjgB6co1uXKx56kIyi6xP/ZKpWC8UU8tCMZIXc404P1EWLIIo4YzFD
uJDCSvpPyxNWd3WUhJmhw1ve9j6jxi1bIqxvDuO/psmIvb2eidqbuYIpWwAREYOEnWXyTY+5HXm0
ZULw9/rQ6ZcNg6feKRHX1POS74MLen4YxkXauW+f0rfAMEkAqjYyadeCuQtn4IxmHbebanwLsYKg
tGVP3r+hbh+qCx+ZHoXFUtPzePwQBbXD4PMIX1tFSObyPRrhhs8xGl2+bye5nwj35m7wDhXS10L7
RcYdZPFQZmwGPnpaOIYd/JRdMin7E9WTgJXcZNpALgZkPjXUZr4wU+V2ddkVPds5eJC0lPjfx7Bc
I/CZO73TCg9+mWGWw9makRuGJKL9Ux35TR+M6wQ7oMLr6BFF8nUv1dYZpy9niJNas80q65abVGdH
8ZBZ8OSyOxoLFFQG3NmW0uvr/xhMGhJWLboM4WgIxuXiNHSM4mIzPB7bRrihfTEBjQr8nM0BK1js
zv2JqVTCrPkdrm0f6QlF2uGiQZ9flIeskFvZ6ambts0gW9sUgtCeQIPs7pK7JgllQTZ3m6yIxDw6
yOSYZ98DzaIwZaYIWuBdx8tNKiDyR/mQ/DEHo2KYqp4rPLazkyjIkOOHLwPMGy/59R3xjErQVHD+
8WSFvZG6n418K0Pas69s/bgpF1w2SE9WOhmeNQIQsu0FKzNT8bSUxxbU05Dhru0HUF8IhfICWUv8
9IPBQyQAs59AD0EXBRsYBOXcrNyytUKV6dIYpYoWQRkZQXXir6FUDgRh33S1Plv7aVtf3A0n0oyq
6YhBhzv9LisWCtJ6W5tWruEY3HigGsEOELWtDaxPJr40rWgEcozXtzz7+6GiyBia2ZWsSJi12gW9
jMSReIagdvznMsPw5cRsbFsHyWjkLVRglkI73c6+tDNEsfKKBPrNcRLkk444yQ4bp9E8qnV9AC3L
HF6qkllGky4HK1imx/zjJWSHJ0qJ1Tx0XVZD2gn5+8C0xk5r6Pqp4I0puJLGQo+QNGTMMvVBfRrl
cpMJg7Im2VR9nh381GoJP9rzxaofajwc+DxofDjH9lvvTTei1hf352XvEZHg1rMi5FAl3SCrmH12
CYOIOkOrv03j91tSOTuZgjZsnOZ2eg+5ZOAkHb6UQ5ntXE5FMykqfyfPfMTTyb7pbp1d/XTRzlmb
x/+BywkPCMDuIb7H6dYcN//01s87rYpgulVMCgHWNpjw/PF8r9FSs4GgNlZkPRXaGMMB6qDddC5i
RoURTTfXli5j2s6rilb1DrkUoCdiNprjkMKHoR3cPy4n5lkcYjOeOwIBtdsqzzuq3/Kmhl1erjuz
RChVPHy+WkHqxdWtrLXwXuBKiT7Uyrpx3ZBvV1l4JVOWpBEowiQo7hOmj96LybkAGeuegrue5Qiw
a6Cnwyd9xyCX4f0wuKK+VFZfSajMDYNiGgow/+RHf9R1xePVo4Jf1m4Jjogak89bxSYCyR7BcFky
U3JHbXbFyMKuTT0ExE0kTHommhEvqC7pmccwNtHchhMxSq48Dnxway7dGbtoSP9jSm/ba9PwmiJf
Uis1P8L9Gpf5qK/kxncFSNeHN0Cr6FVYFpH4PLctd8bmyF+CoOkSN2/qwD2SOijqfiPlEP/XFLXZ
Llnp5oePnK1geWxoroD952KxFhFFup20PdTYV5YxOGQP0bcpHS/u2JXbe23CPsPqiFiFPSB/hmay
z5hm6soQXf2oBWS++jt2nzi6rDjUBIzG6gXtpntnB1K64CM1cCcAErDtTA4tAF9ebnrzWqLLJe+5
jKztsuwRXcmy0oJPnbL9urHCKRbm8MKbRAHsK5Q57/9/fR3ZFMzT8JFj/UzonWWONQGuYzG3hLAe
5PRn7D3y1J68k9mi2RL2ZzivI8MksnvZxdhNUKrQIPsNz8kgv1WFUtaydylUUEtBfTQYTTS/8qhv
lT/2BMGse8vGk8Y9UbOsHCGBNpnY2MmvEk65rBmQJWmj3kpXHEVt0JsY2CvwQmG9ARuO6Wz2X4zc
Oh3LZPTVEBec8xWG3333FXUf9BJE5i/+IR6arPjCY9W5zbbEpfRplxU0nGgUpGJ3EJSSZ93wLX1S
UMvf4YQI2ugTaw9pUrN8Ue2cZfiRn2tozlvU0sn/TFk8AbrTfwd4+YjZmcFLhhBzX3qaV8dWto7T
tdW57EJyLcQ2R7r5ALjREo5zBJPGFQ8maKvxteHm12lfHCAX9mmFpl4uy+SMPZXa1ux+s9XxAMHy
w6k7OiFXEp+3R+MyOdXbBEhuY/S8rU2vn0HFvF9O4H/pJ0Ix8nVFVaS00I2PXFq0EiUP3W3jP0Hk
H1PoqKAbY5WMpjzG0ikT/vxP5kYTQoTBdermCfEVYjvArcn7ciP+3/BcRzPzgZHwVSWrpRXkhNzu
AbzlQ8matke/NwoEsmDyWvGMvkE5rV1lItT2MvzKJQDTGJbfTWkeG2NYUW5mIMWoRsI6QuDDrEQz
R+FfO2BObZkq9N5x12/l0NlwwFEbT9d9iUgOfaCA1y8q3/vZx9a7+VWV4f6CO0Z/FJs5zirabMDj
pVJGzCjj6+efSpd/eR5ZvQr9u2omm94krV9DMWSMx782/gEww6+CezQd/kay3rY6jCrRA0TlqjZv
OS/fWL/Hqpj+cIDfcZqEwYSqP7yOuWOheO+KzZ0RQ/9xPDPNK9CP+3mrJO1dcisiP4pF0+xknYnr
fM0jV5KtDy4Yl/Vu6bSiKidFUX9ZFMpYJiVCNgPShTWOwf3yjD3MV5RlBm1bJIt5eVa1ReMa/xkU
sKOivzwJ5TbqGdk3rOcYSx3sNYPdszMWaCTLqKbDVcsMLJ8kvN3HySPjZapMqcoaLzrTytHBogZv
wmal5My1pBOiq67VqTqnmIYgDQUxYY+ysRUI1Hm5W6VRJHyO3XDpY2Rux9/Zm8l/ExpRZGTU6leP
XqfAduYIhPGHBmMbuu0qu83qLV8HhUCFhctrrsTPhpZaoyQ03s8pNBvDJQus4O/q0AonXRQ21TRt
nnGD+HjOZ//PvSZ4kqQxfwEvJn3iW70pG3TpBSGOQV5I7NR2oSAGTdJ+hvXOes9bb+kXBBfrBFZ5
6zu+GnBHfC8Zvive1jmmlUjPzGeMcVkQ0UsCnRMIxXCZVdsOrqzHIvvJuGs758nkTwJ4L5Kxd8ON
/E9i8KkK/Dw1XtwkY6bq5zZ3sZjEkgMDLtGKk+Jy/gJ3zH+wFZGyqLZq4VnjG+a3IOBwXqcV6cCX
IUZJntX0814u5gJemQ8t5qzU+Fn3YIgiNuoArAkMGDdd1exouFHlMs2IT2cq+m750vYjeMjQtqUX
0gIdBfKGRln3dvwE2xLdayw5hqTbIZLi2GACX96pDHpICUiIHgkPgcR1vc0Puwj7Nf4FOGapP8j5
0eKx9yN7YJHi7RlaKZQpgU4/br+Anf1n5vMhVnH+vfzJYlnntw5aEhUZeP9lUDv6WVi2LZcsWzJ5
yh+i4Z9asSX8/AJQMqRQ1n5xieyy2cOMqtOlaMKX47o1m0OMClkPvSkEAV/eNlet1hbXAo8MV/sr
LRfx45IiWDmBPX7BgTpx9x6h3hp5gwXyYZI90U0Wp4+eo/DHvVmfIlgf8gEC68syQ94G+AzYAT0i
W8NwTeYOyKvAgUUpriBnsm7x/H60/byrg5bwXdDQbhquv8XPsbpRBO/Q5GkJk9po+OBZmOXYuthi
2vs7J/JUHbRO69Samuxhqub2EpjNMzT5ilDjb9MAlF9H7kEeK5xcsYMmhnb8y6ExI0yioNoGJ0Wb
+zWVLJPYPSN3Z1lXPSEiY2Lz3pbHMxf6FJs4dWDDFTGDdfa0ROw7IhpgZis8Z/4rRaS7oNe0/G7E
phDvTfvlJuvaVqIWIwdBZmC0t1mILFNwKXZC2bvoJ0RV/gnEwXBTg+YxNyB9VrkvQzhEeQnBeVsc
L+QxqnjRgnfdDl6n+VBOL6coqra10E+MJCLz0zrmqEnBbbSt/pd1G+M4YqkOmwTS6LAiJmp7Chby
YnYwnMyuevgYh8shQKKR+beiEkEFMDMTpKrdEnyfu/ssYPmcUA+kpWRQiBtbiJcDM2c1aJDUDNiB
Caym2i4DYffOD03ZXyLgiTOmKe9PZ9f5JAN/l4sbOMfu5gihhqQ+pY20DrbSkyMRjZ7Yh5VL/sqv
UrglP6HGqbvVDa7IgSzf5ofxa1dZVCDsmIwV2On1IhDp+Grt/dkWRn++FY2Oc7mMsGMcUSsfuXEc
9R8ElFBs7lwVMhh9AbQu6JoEtiacyAic1+oC7xr4P0p5PiTTsYeS8ri+oHVlfLPKxec2yEUXOIGs
3saV3f4s0i3yp3d114BrUxNCdCZxR55lGjGTGkjZJ6lqa6lqMdYxBtNZ+9zmOzgxvLDqrCl0NQ4y
6Pe9MZTs67J4VhzIirkgSnzVUThKowSMe3NSZS4fp40AOBiCXF/q4iS21Nwbsl3SInlfPnK15cFi
HwpZyihP2Mp6/dikNoLF7uCkyJJXbukF6Nk5bzrQ7ELLdhnM/0ggqiWoxKr0Eyx87HllaBgCVTsH
Bdo/6tRXcUbXE3FQGLgegQR/M/szP0vz6KxaPc5L5c3AVPw+O3Eo3Cy5syESlXlnwmS2pnaDCsDF
rkRw1u+u+7jWj+FRWj83tvWcVOkYsJdHWk/XsiPUc03zACU54W49PeYgQw8gz/piRXgkTRQezsvl
jWgkRUsAKtVpv0OQ4gi+dPQEuUiJggp0RF9wfcqO9JwJlWxADBVaPv4Odu7PuZGy7EECkajoLseh
CWfj4h+PPpQsUDvzpsg2pIqViFaUnK4fi+jvEmIkwylObO4H+Oo2mubFH76anB/HEkURA1tGM12s
H8m/uaFVJLJpx20hi58Y7BzS00JVw2WrVt0HqUbaWY+u0Yw4+xCDZeLf9CVpHkHK+MrR0YfJB9ab
+sJ/XLB5AdgR+WIZIdUzsRFNLnJD7eU3owGXS/WXpMbRV9N/fRUVHetw3D2eCR0nnLdWn67PYupw
BDhCKbNpYP3tcmxpxF3RNFxNnJWloyOQspXKYcgEFLpU79nO+0cy/cq6Tgl01pzRM8o0f9BfeBnh
HD2ad9l2MfeWC0ZCoJ5zN1ufqgeLaof6bcS6qb6AAMO2y5fgB5iCF0Bsweu4pgtfL141oaHR9sDY
4v4oQHaJTH+PJ7o+jDddKmYLSOi57Q1KQdmPlR2EkVCmFUyRHDc0YidP9sV9wU5pEICWxgjmvoPO
rR8C8SxsD4KJHx8UkeciqgY/YRwoRe5oYkEt5zd22puPllQE9oMpwN+Bm8FhzexBGL6lUD8Wm+dL
G9I+Buyy9yxLtR80WaU0HclyrfBvP6seQRAxVm0MSevZ/wpRvpWLfy3YVcoPMZ7hbSQ+OwvjifdI
R+EsYfvSTGS5IEULo9JDumVqtgUVsHohNKRUMcv8wZFshDaHciGzxlPT0oK1mFBFONaQOsgq92q4
YMQ5zl+iQO7VzmykAjelAZA3gD6d40kzCrGMiPlXhj5OFVMDNZDyhisKEiia2kVw1CrXh3rlXm8b
3npIB2Tgn+FX8AVhF7+tFfxHWunIpceW46AppeDCcHBMNy32sSZ4JW3nRO8A6O7sDJVREQch4OkY
fdSu0sRi8u6UftzDhMv8Sa3BQt+oHKDIUGDrJPGhLe6vSwEqgtxIqCxAxhGdaQ4qpyhRV0bBVfZ9
JD7L7l3GkFnayAQkNdzhkp7n6wHG3jQNt1BPGmV4DX9GTC71XZRja/jLIQJQ0CvE38Oe4ALKDF4C
RZ/dvbY9xjVOjn0gh+lZ4jjjqXD6bUajxMj+pBrdFbE+6ly+w4eIrNId7C/LINvBJRjx83U7f82+
e3YPwukYbjrZkdsp4P16BkGKGrOBzAcuM8olaMxskDvxnySLS+6MjBol46N8h1RrSXwLJZD1gQDU
6XQO4dceGCNZyI9kQ7m+kZoeNYSazCXUL3+0nbOLSeLy3FvKPD51ZPBfg7fPGQ0dnKalT36QjflG
AFGnyv6uDUegK63aFnMBfjJzbDC3JfwPifkcSmlra9y1MQi8hPw2Gg3c0RYsp8W92cbTJe9xhW0t
i0dyKMdRQKdoUHjvPfizb/Fi7AcU8FImInOF8ayaeaKtsTg4QUSwKhW/dRM8/RZQ1YtuVQwUxYvy
VKZ3F80QS4sWPGXkd4N8OED4nAy6j0jBxaTrJVAd5VAsoTy9t86JXyJMzx8ArraSIhR3AeWseXtc
qloZmvcAsrjpuB7Dn+TWgMgb/kCw0vxKkzZ7Vm8lX9tmZ6rvx/jxCo9lh4kfC4RcYucD7aLbZKMm
T+gPQSfFWiVTOOXw6AuBY7PPJJzGvhAAdmv7h5DG5vTHhAHWcDUdMLZ8hIU8Q8UQNbvvz312T7K6
ypVeYl0j41osNdOeTFfi2Dakd2tXM1IVx5xSsdFjZBiRYLsZyPZ4I0sCikt6n/JzczEu1RZLNrbY
yjKh1ZQ5a14vxtK2VmUuFUQgpCDZoK/oLSwJ/Znk/qY5qBWqvTw/CIKmGD+QBEK+Y9Y4ALLV/pfu
mNcmphFlgaiXJlH7j8R1aFnwhz4q0vjxoJhVNL/W/bpJe4z3IzE0bMQiJEc1mZBxt0XaTpc9ibGG
w09nBGIvWP1imdmzlgmgooDRSbPpm6dv9nlqClHLg3WspW/hvpdNsOlmQFGQoodUWQa/aPVHtktj
LoNkxbaK9rttFj6hqR14k1z6LgYdjOrWHJfqp+Vegm8NEPcp3KmADNaYkd9q+i0sLoCiBywuKs//
j085cuJhJtywzIbS1BU4YuIqVuZfhDuK6LDeO6OMktHnQkLVQ9jaaSkKI9fadpktLrpX5T0LPztV
PBLpvARlVJwlXWRAD/ZZfSYJ9rZGB8KcGEfw3GJ4m176OHdKHrqRj+97GGKTvH8nvXt+C3+xGHpM
O0/JJuLF6HXCluplwVJAD8KgARGn2DH2Zd+ZmpIWo8Iy4lm/nuhEq28chrLZrWlo4eqMRsDdp4gc
b+05ZNFlvSviwmJs0KAja8BN2dAOtjX5iOdEPAQknwOdYffPWLTOVt/D300lMDVc8fYPSnwbWMrt
LsnwAqgEpxq2afI02KmPSkQHSsXDm1EhahgJaD8ZBAclgZ7lb6eer9XW6qA9sf3/PIEVYFAFQsbD
X848NatL0hI6QtxcFw3Ci/uPaLc1OkKE8ACS0UrLoNtYQc9yzwP+BNQO4IMdlWMIeISv2f2GwMP9
4ruEBWSQAmLrqWxxb3A3DdGui+GfhGcy2gq/FI339bv+jsvgjxtcMjO54kCz3d9IoMOdUQ/MUxX/
Ol31EOomqlt40EDPdnt5t8EMlWDVirMPCm17A+IL7Sd2xLAXyda70qMtGMqDNMHX2QFhD6itI8Pk
ajN0hyKq/6GC26UrD8PaclmJfucdk4JMIYQskZglGn/Fn5rYrbbqZXlY5YgOp15fp1ATauuWYUia
emj1l/O1EKHDqgUkcanEb5vqCjqIlnGhr79PDw+3fdW9ej8LTshlcxfO1ep9ka7SbXyrsK278PB4
i8OqJGBcs3tn7SQXrTwNaAqbK+kQwdLQ+TCSywjSsH1mjpG8ri/VqIPRi2LJEV8Gq8AeYaxH/41M
Z24GxBWti5h3lnLMQsHB12eK9YgCWPmO7lklefVF3OxWplkjjWJo1tYQ0yXqt1TXyb5dBYpM+AAZ
6Pq0Y3rWexMFGCr2ubnRAx6Cw/DAJdRqsIu2Lndl10TxIW5byuSfj6GYJ5PTCS8mxI4itZlsrole
lK9PULkqv2VYG5d7mi3jQ6SGCoQ02OflkEi5la9bTiFnrJiuSTFmMeteqDfinMzUuAZ9N+blmQOs
MDzMvdSDTHZZPz9qaafAqyDNWmBmMs/jz1Dgvq7LlWjxW6O9s20wamRUY3RHqTtx/ssQjl/X74mE
xiotF6NyZn+g88q4lauYrpAjOX/aMULtgdHxtpfWBahVv1Bl0E4O5RRdOgfKSPN0TjUe/E8sXCqM
H7a9Srqn6P2Qw476vUaFb0+eaJrHm95QFTASc74aj1vl6h4pYsGgMzD6Ox16TpxVcmtgQackiAqR
Fr/hAatPpaCS0f7wMFXvaAPQul1aTCZ6+2hUeV18D1mdBboUGRLhd3RG+qLAehrE/FjymTbfgZwR
6O1ikqlUkktJXQYklifEBUU4Pxzwq+RqTV1KeN/hHgdxFq2K+Z3DYJerUqQOaMIg5Cdfdmz+bhK9
WvEValkzcINwmeHHJiLSVgidmuKjtYdRjjcA29/KdqbULhsYIbXS3P0WX/roRqXgEMbVPgz9DAaE
YPmg5WzmuNxY4TNRcjM6/imxjoa1AF+USRHKUnJKiaivJ6u0xxFbacZkQyJmrPu8Ock5kRnYcIc4
rBdAf/t8NhOKPzpkMEaLURYYvniq4ozaczXrPErSqjwZi7/bDG3kQUHXdTsxEpzfxX4lNS8wXoEJ
c0CKCJ8iZnWn2y/MDNs28Tc+cAK38awUm56afkd6wAE2PdNY2zFFZPxmAW2+534tLhW+hI4326EE
aOyOwKKfM+kn4jwB4BhQnUVIVzJCA8Ivs8wPir2uLR+EC38BL01useE1RMdAFMUPV81I7BXhR75/
jX6j+nww5ns+yhMjD7p4r+lu44ef8rUJRqwejI6liWCfUOOZF1/93+rj8IxZft9MMbBMreO2wIA+
hFnfR3gtXrKxxquMnEaX2OAK/+IDkHiddVGqN+OJT6IHTFfWPGiMfCuQ9UrnPtctUJR8G29QCmoe
qSCX1xtVT51hk6px0ImizbOjSkFzLZDIeUTjSwTucT4S9S205dEJj34UnsyANt8a44bVrgV/nWYT
aCkn+q91HjwzyBzz9KJSFHHPqZPhsT889J15sPte8O1YH64fS2IugT+Z40ytePdQ5/QYDL7uIh5c
6wGTONhW8zCAWNO+XSI5Du8Tu3G/o0vbHdlxMBh/7cR3iEm8esjMNwUR1lfbtHsIwEa1f0Dr0Ah8
hYO8dJsmft6AZOIb8PDrHunWXXf3pVZdPXzuilk+O7ZRiK3Ag9xLX/vrrBnpKXGXLiNVXnOSwYJj
ZVjYYOrQXrVlUUxA9skBU999nnAfIhTbuxgk9tlk0XHJ6e09GWtBemQ9BzTGCdkKIXhgI8m0fQTL
DTH5FTVjVQ6QgMJ0zbonBoWuLC5YvCNXjHgtu+IsCTm9NODZO9UXSiJCXouCliz989MAkjYnFVNy
Kvww00VBdcmZvf7qqmHcGIgC/TRwi7aibuNCt6+yXplXn0gfBFYhnI+Qiii5IL6QhMUjgAV4JU7z
4qaZtlhCNaCsqR0wgRHr/ZDBtDMCb9ThwNmBd/u7O9E3oSncYWjkhSkUlmOb04NN0vHAnC+VtLVy
yK8G9TMPn1ss78LeknaprdtisM7lp7jPgsq+CWHf8gFZHRjaFw6R3bCwPDzneH/xdsTgoECpyWjU
wT2+de8D52h0eEijJlrSKEb8RWXXFiMx66BNfuqqDZZO5chBCd3akQuNTvlIJIA6gwyealExrXX0
HNEw3O7Pjs/QobEu237mzw4wnF+3KhEcxxxNaB/3JwLDo4Gug+ucDQmkrbIonzzudOLd4SYacU6V
RWASNlmPL90RyqRAwYb84bkdHQaKHEWBJtmEGh+odnpxTzmmgfE/JAV+QJgnj/e5UqAO3xjsKpQh
4uw5+WIOwMDJw/FCIHV9TQ9iFzZLZ2lyfN88bipOJHkWbWTbOx4QM7s04taNZZTsZDBPyL5WCfUr
0eLcY22TgmnKwXTHQFJPnv8aeszte8lL/LgSSH1eKVVTwf+6dWkEYdElAGG/R7/rP4TKDeT70tFj
kEiGHhgaNKKKb/mc64An689qe2HfQP7faoAvJAb00/+MubIPhIGUQML7AmQuiI9VwUgQEoMhYm60
wInXfGX69SLunoLJCE4aQeRNchasMRRsr9hxAgG1R/UJEXHh2XjJgV+a6Wkgb/WIP0flclu+zJEJ
e4artdVci3vo3isNrPKYccC/zARYWvUkgELPAwB1SXEdQVEKsrl/Gsi+r7QpbEaCCLUkjNFWQ02P
VlRyCJXRciX1v2kmwW8w44D4t4UswmNHoEexjnG5soxSBS/Jvi7aU7WxOwVCDVmx8+vzPoU8+JeF
ufGsAnYnPGbKCSIw5nOfxXeXCyKf/cEskH630CoLlsf8QzL5ykyLmgBrgrhy2tg3mXtaPgXxh/xk
oCLpYJgGKhjoNB+cTZRu/AyKmjWIFjJMCTpsILXkVt1iGBoCnJf5UiKRQQlUUMBjDdTy0SNzineF
0gXzZHdXhG2iAsyzaImfwTqCCg0VPP8XOBJw34p0EO/ffuNnC56/yxPP/aepJ2uifhD9noogNuXk
8hd6rqmwpagg5KMMJLNJpIFqyIiwhLkzgE/fnnd6+Gvzn6nfTjF+JfbMCq+FfzzHuUuraFCI+2us
TqRzZzKmGGMold93h0NaPx6mg+i0xfo3Vvd2+CDJyTUG/MqdkXennNX2R0S81XZGbVqVTfW7fEGI
C0Pdmcp7nWKwBcVLml13cM9y9rovLlwuwUl4m3YjOi6F3xqyjQLsU17553aXsNmDKtKg38v8alNy
0LAA7fiG1G7RgTcRBiAMVexLja+Dv6MVfNM6azD2syXFiLBeYgQvK8uDyVXS0BjNWEPA3rFDwtlJ
SWhidIDEPpzemZ6QfIIIRvzbuEqLfHBzLlS0Oi2OHtQSNJiukeSh9L3yXppb9uT5W4Wga4PxryKb
1lXX+vbbX1UOSfLV/sbaky6i+gMEIKSWf3ncY5nHkkI19Ig1GI0g2YHYPHk9pYRST/K+IeUxMNa3
3Dj2YZD9llDokT8X7DdocfYgas65A+OQd1OdFVvOIv8ZtFVtvRaiRfq2t7tsRVmZK1Yp5u++/8ze
MInyo+pUF8Pg6I2GXZTzkkFvPiH6+sI6EqVfOaYXOZOyKth1p/2XlxDkY6tbyJ4RK0jW3HYE9vWm
6JBqJoYPhhykQB4EkVkHTXFZfnzm8rAui+4BPONOBDxLiMczslrSWWPK7J72FUPNFBE3wIRO+2mj
Tf27Vd1czsahimdoMw8bfrEz+pbZknHLBVBnU8A3UFbPplheiaxajEoKgr3xiYp2POzd+HyYeF1Y
sOcZ7Q8l9V4wJ88e7TjSwiy0101TRnPA1C9RSULG7iEi3ng2yFarJE2I4rSkXyTxPTd5QVrhAVk/
iX3S4SIDI6n6BBw5ukTOSM0iTYXepbKGEFXoummU14AoNywQWuDRbrgzxLLYw5oVv/GNMQWNSD7e
P0HIgRvoVVOcuPilbAPlXFW2qjLE/jbILr2Taq3t9t0NVuzVC13Fjkq8v7xLRAS+dzecgudEpGCf
joOkqkd8Ota6R2kawVG1gj0ldz2ZyhmEmUHs2BZ0Z3y9i5SV4lGq14EtvODzEfhhHNXi+KeYruHl
zot87z2w/3MPlTixPxiF0omGiqyylnSuF+l3YmjjazFBFwqrV1o4SZ2yAEBQF17eBrGXf3U2uYbr
Emu/K1TauSJru4+yWQvLHqH80WVilBXmQW+a1OQOw9VqrFixidVfRatRlx5lcFsmT2LH48HkdsJd
ZQTJmrFb7UVzwmbOnw6/QX/pp1RrKkr1m+r24ikra3ABd9sqIFvZ1chxW65IkSVrVdMnRONJH5AB
5ClrNQ9oqXNaYGz7MCq8WdUamqaDNQA9L0lCG/XIw5PslY9i9yzv7p5EcsEUNjrbtkp58yPjZL6A
YEzDCtrlRUgExyTDvRdfi/0ru4cum3pV3718R1fD4GOR3p/GuJ2YdecbLr/jzQyazj17EMsKGXiq
Nqs/Df7XgTZ03X0iHzpmP03vxJ3PireL7oZ2NLqAfSwW7egv12KylHozHiT35c35A/pvVY3q1ghi
XnBiK41xuOpDW6hEgcI+DOldAQstTaee4L3U2kIdpsBRUi/Ex/qCn91E6EgayokfMABBscpJBSqz
yzcCeNUCtL92TkDPv7xbcQYWbHqW1T9HLGNgDUiOOVncScJBwUX97C5CTwgZV6Cxf/sG1q033sSs
oG8oiwd8VznZzLaBQlYRlH9nm0INNMcu9Tnz8ZLxg+KkpOWhzG8b272DqFsaogZmQphYc25M3xzK
Y5NvURufkcd0VTCSqEf1D9dlb1Xk6PLKsi043ZulsfKDssqWYF2Xi8zFfv0SgyGfBHYApRkOxhRI
1ez0n4d4lTFYt2EY2UnsE5cn9ROeeAvEjw+I2TLitfg4FkpzOFkwbCIlHpjzPksjFBmg2qwnbjjI
19i49QHPmqVTb0WlCDTI7Q6eiJF6sLbFhUaR0T/OZkxexpF2wov7eyji4qfgRMiYOauACZtofigh
x79inRwMukHgWji7Nvzp7wwBn8do3OFaW77SVyre0lW8UlV0FwmYM5vDCAZ81v8wt7gSlXMkLHC8
0Sr7XMb1AWEinlV9+a6HI1vZwxtXymdd9GKjwUaBAS5xwRr3tBdR1RDRFWjSjO/UWhlCYNzAZa3y
4p7e9MUWHaEiQKcvEyQvBfatERQgMcDFz4pH8iCveZ7rsqeOeCi2af8cS4+6BDlMtckFCLHWmsze
u/MMXpzI9n+V0rnfUU5AmOu74eOSQtuvYvz+UqLZe41Ye8Z78sgLbynKDnmUesDg+ImD305MiIPK
2xBMRMwmtB92XJXcFNywDh8UQDJBtIeWINYyKRoHry5negaD5HJXOzxl+KHN1sLUksVyIkRe9mdZ
LVnwR9CJ5zC980vWN4ckDeVgdkD5SblSzIGb/R07uumWZWculQUy29fqhxB1URNSuaSTDrNcB7dc
detTKDcT6+7soxmdyzc5JUCXHynA67YULjG32fSAeZN82YSwhIKAW2My7r+zlwao+RaSWdNoqGEV
+11B0OhZ+KEqxSzonaHduobI1CH6VqNX7NoFNwwGp/cf6fLwS4sGG6zE4LSU1xod0zutTzhREE/G
rDlDBA+eiayZdFL/wnZtfqkIhxb2vJTqzqgRWE8VBcuUCUCg2yG3w7LNlHOM2wbxB7/6eHQJ3dYd
N809sCkUezNhG12PUTICkEADdvZTksrwe+rBlzR/cWqL/DzXgMHPuYreMp2CfSPIaoY2YyHMBRA9
uXMlT7SXydXMQqYX+l4zhiDs5Fd/AvvAlwNOgk/eLhLB6Mjary8ScW35HfWQxFTaKt1HGy1MiQas
ssPPEZ8Ylt43FKUHH8XIyaJC3Hmd/dn0I91Ev5KPWFto3jlc/9QsSVkzNjKjxAYZL9Dx2+YjhfvT
NHRsQEhDrxFXeu0IDtoOEt6VhpihYMmYPErQVMmlSEi3xppjkEHqxoeLqtfDjQ31TFKqh4ht+2jI
pAwMQmGqzPzQFQhUbrfnz+FxLQqmDzdduLqsGywu3TUsMiYsNlWLS6oaWGUn9fgKhlWe7Iizovic
HNlO9BqQiB0x/trvtXmHCtPpr7mMZ468+7axCgx+8B3s25QiCkLdvVc5DSTNe526NlmyyQpK9zJk
8EahouPJRLjOSxfrvbMlGcf/3yvTKV9aL612unS1U5ybYsYkwtMLs0mPyJ4CuP4MR44FiQnYJ6Je
eT79QJD+bmHcHuhGb6K7ZYBG3T7Dt9nYMFC2MtWNLWhS9iV8gre6pzFRJAR+Tw4F24yN7xJPFqUA
pBFnEEfv8PsAo2tesK8zmqSU1tZF6HcS0UKXkWa/l6U+HMtJdaE6WK2TWbldSylxB9XMKjdYu8+0
AbAFBy2QudCDig4Fz4bDseUjDGlIcudPl6ps7GUPaxyinyiqsNa6pbzr52C0TNL9wTy7wDbD+9Df
cw8XQ/zYSb7+oqWbGcaQq8+8WjyZgaHZxJr6kKIeNAU9bZ1DgFzYS9AffEWB97D3gTMVz9axFeaj
mAoKnxFyhL+ykKYzjwOA6oIAXbAX353IbV8SVXs3PNG9uwKPc2RBX5xdlVJEb8E2KP05NxXAx6Ji
sjVPzakRHM1gc6siBMhh9OytNz50sLRsguudh7FcGDgTajWHDTxpJxCadWA2HdRVKFsTwYCXTuQS
ZtgcI9fhQEcdcqk4zIZGh60PjwCDcNmuRFUGQHPmgk6d2KC8xI/61OohRInotoPiE1dSLyfpBQvN
ytrwiN9Qv6gD1mtfvHW8ja3DA9owjo1SEN0l1O4OrGETyAOvrBjpRpYL1zdktykMytCCMgHGP7Bl
zDzRAYtntVBMJTnz/LwhIl+E0tsl6YGTqm+VqSspBT74jleDb9P65svWOE3p11CWbowxlndknLdA
ssLWX09LisFYTjEsQeYUbM40paJFGIILhiWMiVDnHaLIqZ87RlQqL/rC3ugj1jOCdPEGE6EkdzgJ
DmWRN53BLEcgdQwxFJRTOzGa207fvFWXc3cTgEsYovqqP1g07GRADPMptpr3dr0f3ORHKo7NyhQQ
KZEZyLiCCCH7cRAhnhPUrQFLlWvI4B/AWdxbL5AK8xzEjU5ojqEaEuicG2dBHY3qnDXNKpV4gyF7
b3E144EtN2N5gSrWC4RveFYI61Esn5I0W0X9bYp3AynCORLtRKy6L/v2gZ9dzDAedkxNWMx7O+q3
BDZTLLe6xepzQDsjbtwKpMa10LgcCLk2rKnYvqVp5sCdzOC3iY4nKWemCgLjgvy2FNb83/jnw+ov
TiF0AVFZJKRRpnaQR3WzpGMJVz7/bfmedmfW6E4Ppi7fbJ2n2ThYXFx8/UIzIEyVoV5SBlhOGJp1
pEtsAii9O3MlwBIcw7WrL5m2fd1TJqhozPkniewBarf1Ng9YcdjS2NdCwI3zXdsBKVBKBDj0Xr6f
bAIg2/KGjHB2c/VC7z9moc7OVkHE3j3ZyLfrirauGYI4UNW+LBK9y5k1YA8TcwyYdKrT9V6SGyRy
f5caP5XW8UEN7eVPsvJVoXQ4bnpLrGpmHr1T+L+jQ+eqz/fGlGnVPIMyNCe5CGqTeL3N1JdDuqh/
2qoKd9UsHIUxSFrZ1p9uKPgWjvGTXArdiePCzz2e9quGExwXy9t5yEZ8c+w6u/uaOmg7dTPj3qlZ
/E5lIPLAgMNFhfVzHengg7PtnHQGWSTioAY2dlbXqaKpLzFdfxtOv/+zuh2D8RhVY41WIPN+CqNm
U1+nSDNGSRHhTdNU+mysZRQENcJ8RzgFo5rbIbce9jdALhle16p3mIkQvzyFvZJ7iqWbP2RxPfWU
I5u5CsVNZoqc2kGISEzBj/2rjSWJtE8ihR0l++ypzEzTvtJ1EL/pr1+GSQkltXcT5o6ZlPqDwxzv
ko94MG9dDvS0rhznPL8doIm+WW9xdHm4VmOZs8zBuQJGOLo0wlVKSBL4j46iM0sfTTadAM98y0rT
9O3jgoXAM4RY0UJmNvzG4rXHfpdl0iQcAcX/6eGdPM6smx5LPGwyCwdsNOeux803XoFVM25euIC0
a16ZVRbIC1zzfNwS7z0rRRtV8iAZs39POMSVDZ+KnS4LXMQw5ur7ViA/Eq8HD4Oj9hUzOU/uZOqJ
2RcmpBL7zAiyad1kFoRWrXkvmQOpzf3lUoEw12pyW7nxek6EsglLLS3VibuAwi0PXjXUARCn7qEf
NYZPWFKhVmCgEALahLGYkegR+u1M2TIt/gNaIRhtwEBlYdNnmsLqgyF2DQzMagoh5i50pxq+nkBd
d1UEpJIEQT5RoSjgHTEi4CQNiZjLLshPI8HGZx8k5KenZ8RAN8nqFUuIFB7BrLQ8N5wDgERmwg05
TI7NP2+4nfmfR2PBl/lisIx4gJHb3M0Dq7AP67Agj58pZ2Ye4wpgjiHc/rCwOQ+oJG40VXEsDW32
TWCcQKmuEgzYwxydmf43UC73cOG6IVW3LC7VaBtDFymczGc4fGNgJQmqnRN4bs4+m3+0MSq8x7Fa
j1Fz0XL9czbvkaKLVNDWOkaskEKxS7yxqx8/Md08XNB3r7O7lLoveMsf3kenArVukX5pQiGvBu9W
Sf9dK6yCQOJujaFhnlxTofJbw2Cg+Rxjk38eRswTvbrhU28zKG8/rY9PTa2MgeZC36ceWLbhuydI
1rtmvClv07P7SYu7vwlusX9sF+R0WA9pfo/mMI1CbRJ2KY2xzo4xswzH1EO3gBExma3pbetfYl5l
cEyjMqF1ZJMuWjka+RPADmBq6XLtuCF222VpUgfGtdCtMIFuaP+vcY0M+HJB59hgDJSBZ209KgzY
kQxb2p4KUHap5v2aWODehPD8mBcyViMT4w34Whmsq1SDVzRdJD7We9/Vl+tuyI7a10ozcueUCvNU
WcNpVwkPRAh1k6zOHGWhNB8LrDzpu3w5dYetMAS3PmJyQBEBEGKaEJlPlVAbfQs57e5glEttSWsO
QGmLeaDjyo/LhF91lklFhOsH9FVbo6xPCv/rUw6tiJu81XPy/OXf0rBGuA+nyMcjJ8AGLV1Uwlcw
0ixzmw3a8BNKUhhMZLH/DZ227jk9nQrSehWBOKqDWnLdtjYWHGPZ7xh5hhVGMIWorR1/6YqHE+Fy
7jyuiUWfCIvnEcTf6zmKrVoB0wIxvcRzz8d41L3LEmSYfaVivFBpIMf/UACvWg6ljxfxCDN0n7I3
5+vj2gWLEMX7HSbOZWoefKzEqQbFN9i4eSYnDou1+XFR95ErSbvaC0v5mWW+/EN4fNxUV1/bvCPx
BzKmueiuYFxrgD4z/Lv+2YMMj24QrmUlCeFo7ZudcSAvtfBj40htO7wzQdORv/G3EYsVFSPX/mLt
V7H4uocd2I4WbPJJYbj9XNqUj53Z/5tS0ntKglQHqXvpeiZsBP8HUtX5jp1WNCkIibMDfE+Nckfu
npbn7Y27NZA6YUWx8/fwr4/zdBxccFAm9zOQtdlSVqpJaVmDiSDkl5+0PjZYBhpGkpFo4DqG0P7c
5u5Ydx+6K7VBIsNrdYA25PjlJ2/zNxcJGcukTRbhm92wGCDhRVok/pYHmLfOg9mhNqsXaZo4aEUM
lSF9BGoVhZxiw/uOWwAshliAdTox/JT/LQssHEf0vLE6pQj/e0yPHgfk3lF+Rv468BFGa+gE6peY
NmmeWzbXOChajsr2iTANdwGRgaKUW/z01fkB5mjIFmSI26uGvzCmzHwVsZcsrUSBAFkZtm+X8+Hv
uIWDFYdPP4ayyTauYkRIvcP3qc1B63CAt1DTAQRD8Rwn+Gnk9GR8Jx/LD0CIGvDgTpb8LhclIIPa
/FBbV0pEWx5TBPM39DzTRRfpLe+emo7IfhJGLDLDgLJckGwNjIlacSrCem3joIVSeC+tsIwkdBYK
E3BRIi1DhpihGLJKVeTU66jYhfwbAya9jzs8QDBkMZUqAThXCgxYj1hzY4ld7V0dfJS7ScymGq9L
KDkDx+BoyMHO85y7/YTtDhtcBxn3z8RhatSe7JlJwpYd9rxcyN4i1wD4kFDeFMPTndpCHpDNpoiL
zMS9hw9yNT8j2KbjJRmPDzVE57J2VtMF8tehT7mI6PFK4D7dVts9joOam6Q5h8sb4fcYTaVs5dgn
81dGjN/VO0D1Ly9Ck3NvcqC3z2uigsfj0A1QDDnilqFE4pM8SFYoi+Jc9cPxxkOTTP0ck2te7qK1
vJMlxihcZmsOFOT5Bua/V0evZgNn/ceBTG9IyEm04spCQcYFa44DegOK+Pct0hIU/6QCs8p6ggBM
H+KoKSkvcFSbO9t4korK5fkVVs9oaFh2Kqx7Sk4VRLp15GXBGsnkwECAvXpfX14BAsZBKlYGnvYq
Zg4u40CRjQSQF/INnr1mPvr6FB/valSc4QvJM5T9cgs6KqeuujGRDr6SVTca1mylx2Xjw+u8IogS
jw3kcoF4heYW9DufCPjW0ssdI9Q5xskFbRKEw3aPqIGLrdI+YXTaSypcUDLv9X0MhuG0sqvSl6F8
8J3r5R5VGBRvWZvZXD3J94uXHFmvdNa7DPs3PZi40Efd5PpS6fvuQPn3UiF5oxohplLjaxNqaiP1
WRSPB1qsgZiLacig8gT4vSaXIg+DzT9SGWDkwNm5EwRTHdNaPcbShsNk2obbJr4YVQI0Bgnl8FVo
FN7Co4ln0Cs7xuOr1mztuuvQZpcLqXUHdO2PYB3jiHCRBKbfKQ3QEmLPHQSsSmL1qJ/uigGQgTt/
22Glmv7sRZMPkiTHqhTvoLDioKgAbrXHwjUtcJ8yKLUhNUa2/n2w2c/7Kkstp8ZmHvdvAZeJV/Cb
5+7/kdFSD3U3XXe5rDn7sump7QVUp+FSTjfQLRhfo/cwUm5RKPlmQ2hawYk1R5V2BfFXI89g15i5
yJPzBDpKdkri6Xs1XiPXM/YeM48mve+tP0eRmL79ttEpuwyyHJHoR8DswJ7I4vfwboGXHJwOVnVi
zV+W9U52SPt3nug/qD4flkX3bQy1m2ssk6n0xwPwhuqkpc62q3W4OXN7Zgg0kBkx3m7Oro4R00qF
jWUOk4wSefCcSa39QLIBW8XubilUaarPgNreBpz6eC8Odjcb8V+QJ2jo0SD3lpGrykJwDC96rrk6
DXhMjnropfYN6+0+DjF5f2Lt3+sXCsX8ckG+O8e5HzUMoLMoPbg+WjpJo++3zffBZsfStVZcLj1A
pIAZwgZpBP39cPtFcm5bgzGbWnh5gkokHwlqwYogGvwYgYyeu0o65Eq8UsOlrXcJMEZoAS+iJ89L
plCNAK307HtMDyZUNFDaRHzNYIrc7fk7QhUAbrBFX8RmhwA1o3iGPAJZ+Pzl0ZIvEJ+C7DmEBqpd
Mu0ciJ+rbCY0xbcqt9SWuHZVclXEU/mg+umJlHwcdZPs99rCXb/K3unh28USl0KeDJ2Qmwz2Tx1h
IP8+Ah1rAXGZ9RonTokJSa5KIByRFNC74hvKC0mcS+9U+y1ExAJnCE7jPVyyKgfFXio72NsdMHjj
wxxQRkxt6hG5FRFs5eaKXo6uKBoEthJfCMj1G9MTTMsR0kzy9NDDdkyFKdlVssOG5vQr/mbE+SVc
huMcwENkN4ldF2fsNpgaDApa29NbJEc0TSl6wld3bWx2uJ0EveZ7q93pq4SmIThbFSUfI3C2j4F+
Z91Xfjh6mV/2AGDkSpkoMx5z3zWjT5hQgPNt0mZMdkkho0+0WBVSYk1iXszEF7mKhE8OE91It8Fe
Fre3MJjhuMNW9DOigtm4xiuzGeICSiayqSuMstnaYJRJ7VEhkLqKogHflU0sUi3eX/mRwdtdsQEG
yDtOzTbjwBLZjqieOPW6YHKeIjvKMGs4Fe3NKCJnS07iJjvGQcXVjNBJhlGNkdt8wmm8zluaBESq
QlvVZU3hDxbgMbVCESOdii8w/jDDl8QSuHzwdQQLjbHozQkfhdj71dJv6Qj4+Y0xY3993W6BeSzS
cSS+kaY/WEv63/0D9SYRNxtjnU8di9DgPiXXx+4fA4+LS8LOGcVZXPj0lUw4LZI8Bnb3PTmmb1SN
jatHLg7zBK5fQKYMVHpDtrnBeT+K+a7zI+n0uVxgK3Wu783L2x6R2SajuVCcmteyBbplIghruiVZ
3K33tbRrK3g8QsopbEZWY9VnOZMPRoyD+owZKW0grWu33ZQh5VS7y3wnZWW2qR6kbqFKyTkfRzKX
zjmCQEHZ/esISVqpR+pgd1eDZZku6ec+3CCZHPzD3o42nd4V/ev2WjyoteHEX9PQ940UUA7Rufwd
CHrhQAKtS7GS6skbEG6q7/uSdkhBAZ3tTNcsw9R0qrzPen77/RgsbOnq6Aweb/Z/CMIOiEE0vUdR
uGjx6i7ZF1J9QMbPGZsRchwHfiCT7Tb7RHmRJxePWwNP4QKJJ+nu7Be38DzNLwUx8k859oPrxKOZ
whmjGaWRFAVioSRhWIxN5fF3nSkg0RRaK2MCZR9FMewbimwk7hOF5dg6VaIN4IYZATOIamJh4EMK
xqqqaCaYPjyeZn1TUy2ps1RtEeqnvLFL10M7KEcsvrPaCTM0eTyCucSFESPPsw1gCiXnUBYINxGL
IZ0+SGHMULuVFB6ZTbXjGzicx+G75+umWnaSgUas8yLixqyXe5Xrcrni26U683mdTuuca2zcyByR
Sstu0hQe8rY4aBhjx/xmlnc+yi/qc0gLqlO0RvHFMmKDBY3Av6t5ltN+j1xzv3AVXDZOW3EMkXpb
xWzB5VbfsQ4Hn4RHNeinajBPV7RmA/kntUEKlVRWl8y0oz1caKp7ZWEUus9sxLfNgTszDRQsrHWx
A0ck0d96BLA+cyuXxb107SNKktij86lIvSRwXmuH0BY/atBFPWaKyYH9QwqsoykwLNZhPy1kYITp
dG+do0GGNSB3At114OpcgmzodIUsQsITG3BsyMk0dbtPHaZnTBAZdnvE/pDVIeDAF7ZH1Zj7KTOj
aX3GV2z7wX8n022i0PjDgaWZW0OSuYyOytLzuhEjlSCdgFqoEnSiIZkbJL1fpz+f9x/XIewNMGnv
BkrSYmVwh5IVa0T3CA2B8gr60qCNRkHle2cIajPoIngU2Ywn1ZSmFpH+T+wpidPtKx6iymILZ2VW
CR7j9DVsLUC+c5q4wQwlW1Y29iyy8d6+A3O7WalFQ8uT9o8rpH8JYQhcaY3Jj76L+4QLL8znlxet
Zy1T+nvOtUCh8ZmMzmukD5EwujpbhIS7iJLxUdap8xHvDfEZrDE4DDJ7Uu/AhA3vjn02QIndA5AN
1+cQXQkhyydX3/XihZ+rb/55Wf1qt69eII0xSNxKC2mdPYdLHawyjgsqpM5DyAHb9rezUAMAQVZO
HqTTuSpTRfu9pK5SZTjf8c1Nm+nxq1wUyqmlxtcAf0gJ1ZJF1xQkWNVixwdBZk0mzdJSoYk6dNlw
YKbIPKIEmSBI5sQtHMaThG/HSDd/W5XKb+Ql+Ejq2APsw0a/SBtNrPsUsdG8YBBOXsmEKIHTimDU
XhcQuKL7UEdoL4Pi2QymTpiCsbs+LrZPOSAZE23+PtggpCUdM2IUocovseUcToWF8QuQrCsDVfij
yjo3nNrsR+aw5eerjbdHz9dTAERksbB/gS5NjZNIa71y8By2Jl490E72HGfh/XfipnsIHmoh6MBy
JxwMCid3C0izHXSYyeqDPRjmhtEZVN8k7/Wl91J3ZmKiPzduExF2G5DxqjA94+EUK4pG5dJ5Rd4R
PcCeBLuazFexA2TYKyWfpsEr5SJafiUwof8kTnj9bNrF8qN8Ycr4sxc3+2hINlat3FUhEpGrGKIj
e4gIa7fmsKeu41NfYVeo+8qA8gJ2itGjahi9u7lpiV91NJCxYmTWE/wkOR1wfCocqvlSc68GA/Om
e2UvwR1H7+XQ4bxJgoTWLmbOofbH6KYtC9I4VSg4fvvVlfpRWwbY5gc6MnJNybBktIa/T6nTz6kd
zLbWZNe14vuSI1/60owNAQ6Z2fnQpYosxebVGe4+HFC0hijVN8aQAAi+8uq3bLT4ltz9CBM23SSP
KXo3fSZCfx955fqEJwJG5E2gTdIOuYh1Tic0cVd0tGfRo6A4HhjEr0XtfJPdWqiBKKRqDuhnPmD0
nhUuiYit7chSd9R+iBsfmDWcxGd+2eq8Vr3R8Y4E2ytxI3uhUKnUCL0r5D5rSn9P+MZ7H/0y9zFr
V7ILM4yVZHfRuyVQHjaYzFeXNiIfiBvZmcQJTEYnbzCrQAs1fRqQt1bKHOx+D/e6DKy1DszVi0GG
6SJ/owZNL7K5ADgZ36abEpTBQ+rs0eQSsUOo1J3aBK5CUz31DWvXYMs2tz665qMghQVVAtRiFebD
bHLXRcDdQJe1VKjPxy1JICxJbBexv3kvPSKgXjX0uOpPfjoCW05k18YyqTp68U+ERGXRwDcZO6p3
l2AanFRn2/uqxwLd78vJbsMtyo6CZ0TAvIaZYC7kajx6Gba1V0R3VTNA8/3SMAzYJWivWpEm6g5p
AbcuIIqvM2FPRp+Y4H4FnADczPiYE/sKhsrDKycbM1t6A/aDf+CqWW3PDExAtwRDrLjXfIpQnXTq
oApXA34UVV4jBrnjHn40P50Hu92NHs7snQOEHHxZbV03wneUOhINNh8ks0ZYwYKAyQJIaxXGCXOY
h21TNaLXVs3K1rGlq3EhneNZCiViT6eLo8YuEiIixZZC7gnpL2yxhx9YXv6uj7TcZ2jlF99l/Eyv
wzqzatIZ0u4fo84L1Qo1qaM59P0WwlT3IBCHK6KnK7Qh2zzkW/yZa5p6pisvTPktHYUmt+R8RWYQ
YN1KTpe0jrjwceoZkxkPlBPio/yLcayelc77i85Obe8ASX+xVoQGznLbXq/BeKvKnmHvW9Zv9gdQ
JNdADEP3Ue1bEugdKtW53uWc36gpABxaf8U8CsRky/vNel+1+njFUEDAZPJRzyVzIF6NC/xIKOCd
tkzN6TihDgnoLnUBxamvWpBfy3nrpSYF7BvCQexqiiV0CMzm0jG29rnQn70bwpBBlRv1E5fvjHyp
zBxDhXPZwHl/swqY/iAA4GfZwStgopApOo9ltGzXOiskDAwGmNlRIk0pL89Irm4TiVUE56mWwYHO
2q1dm1ZM4KykqaCpzQwQOp2urgGQ2BJNNzi0hutdYs4o9Yz5DxpSmWgQXaXRgMviXCMKt+oYGBH3
Bm2lo+4F+uuAPzsWzkzdnX9/Dg6hukfh1Tu1KewpoPv1YK+NpZ5Cy1JM7DiWMX+ZAH1o2Dn80Mxa
HLrxxHSQehEz3peDkSpCPR2hCGSwkfHmRYWLRb+18nUXHRALxIT4BGube781qZi+pzmZQCD8RAvC
LrmWY5Hp2+Oi0VmVgcAwDExJrMXSTNEGBdt07fG8hCGUyG7bWN47k0HjnKIZaq9JzNLT9DHu0xAC
EGlMcQc2xP8ZEdFdAde/h123/nKhHn95gC+/TR3QcWTEKAaJ/cAL9w932KR9Zo1WCrbZTABHwdM4
vmKecAa9BSwEr0ltu4Z1SQGV5NqPQVfUMZaADUv9Z2vbSZi5YP/fqtTNpDK34k3bB2qGL6AL8Us1
2NG5QMd2UTG0QyzalNr6sxseCx373VCQRlN/UBiiR+5JxHfCcNW3KIRhVvujRM1f7yw0+SnzWegC
ABRVAOKmG8hp+MRsd4xNFZz6gkvXFZmerVZgu3AbRpupgde5SF4Q3lMFFiq/xJschClr1Gh+NdCY
ZsnSIo2wqMIt6cgMfkwcOpWCptn6T4WRFTmkw8FUd+Uke6xNEmzvD4AIkDNBh0AewyQCLMIP6oiB
vyAfpsfjaLdTS5Ggmz8I6bOqAzxxYp6JHp5xiHfWu3Xqfsmk47wB6BcFbP8nHlwpr38I+aEP/9ki
ZML3IyhgLg6uf/H7tDdY4LDgcPqTugWQEF7d8b9o5Tmod/bUjF6IOmfi6/7wh/KrH5hWQkf8G0WI
aBlCZAlCIlBlVf+KrmVrSYrsZwMV6qq9YojrYG88qoRzKa0/QxMAIK3GLKISLDhcP0ZOuvf3gtVq
SYdWpsOZ2q3izWxJq9v8T1k11tN1FQ3HfNpc6+eTozAHhwURTWNSUOL5WXwge48Ce5r+7Il+hQad
IZ9oH4kmiA3k1h+jczijlCFFv8OWtejJO6R3lnrOlmXVn2DnlVj2I9uCPfK8IkOoJJOszMZhj9a1
M7dZ8kWY7K1qchzflCLMw07Sc8Hm4Xo3gA8fV6ry/Gp+MJOGR/Q6b429RvTBo1Hrcjs5fJtyHSX6
mtZfBQyOzA/384Gku8D7v2NBGQOfQBC4pcUuILwzn9fhHLUnN61Dx4mfBMGjINPJd7/asMbxxmcj
lPtjQB4V2u45R6QN7WkMPVF2R/58k05IS48dvYxHulD6EDRQw6Zyy9JJQX1p0dV/83z0arrzxn4G
PtZ+gngpJL+RGeOypPnj3iopKH9AGh0rF3EyO30QwMe1/fOg6mHawPzRghdGhh/qeVy2zQRsrG5y
xA7xbPlicoAsmqbvvMhv6J7iUIBaemjKLH18wpquADL9DY0yMBNY/Vz17JVr6jn4chWJvo2qzohQ
1nGZr5DaB68LpK8YMZfN5a7pvzOxNpGlX++JU55iLkcNHF42woIkTPgXCWJ4h67pfJieaYl/yDBj
IVRgOzBmDfNh6+E3A3w6BVQngCpfk+NQ2fLacbYuiHtIh0n/dOX4lW0bxskgfGIQd0bwAJCelNc6
NIr3CIfnRxLHWLdEMKO7X9lBUda2TObYDM6DXoIM1g+R8qQXKQGsXZgAlt8JyVVbiN9Dz8E4yqHg
QiRPZVt5bE3KbLTD/zwScXA2eJJjCbDiyFhOI0PMss7zi1m8WSyjFnd0HE15epM9IL0o5O9tBKrK
mycCyIfM07yTEHKhAT2iFXsHtFVM7xtSpXlkoLK50WXwvs1SL5sCW7IqAkJ2Plk3PvEjWf7losS4
/16Ok2AulsxPvFUYFsEttlKgPYrgo2XD53h3bJYr5kxUIoE+IWcxRKkW0fmKb6RY1OZqxIagWMKW
P3EjAsbrKam4CcSFjBQMFMSAR/rGBy413+ifb5fEBpI2O+Qd0HQeulG9OD13q4Y/PsUz/V8xsKS2
qcMGY4hmTJbUDT+J1q/jEvxo3m4T+XGz07PjVvFDdv3c+lOh1614a0FYiPp5XPkyh9Qb+N18pvzW
yxl4jUbgNhEK+jshjJQa7RykSfyhUGJrbKK3ehmvqWdw3K0NfZCy31hYq0wk6zZ0I5HzC3ERkVhN
Ll8epJQu07E4uRayunzbjBtcqNoo47zYrUBWAKKT6mTxWPW7TdrROrcolTZ9IkyRKvDZT2kx/Fyv
0J8HajZxeovG6nB3gilyxPTsRjOQlavyOXC8vn9gi7FwGxNp4qTreQ/fGWUjhA+Ocyo4MAd30DxY
1uO7o+fWBCQpBycs8/LnrHxB0iOf8+/IclzTT7hQKW6xMYhkBWIUZTogFrSrZEEjRDPIpWkYq4Ns
cxL99KfplG+IDmwgGPQruVydYoSQnXhec5gkUlnA5zQSAxt9tJk/MlCQr8U42rfalLvmYTTfSf8j
5mIkRZEpTbs+OKXnJNd0hxlvkijondAO9F/PYoA/9aO3MWzz9gcx9akbqrZthmsu7vURo7C/oMlf
AYAXy0FVAeacQQ7N1nLZfllgQDHNy2MlMEJNpJl8bOM5i/6Dzsuba12+AdPtvG9KxceV8AbLs9yg
A9o1WUPMTZh/0HyaYQz+px2Pg6lmEuwEQV8dsfbnWE2V0HQavetNITY+tVyo+DZoWX2ZTr8No7al
aODnIUmfQ1zqVtSzJcX5L5RSxUe7o1dlu5yHhyh5n8/iEcsBz9JhTEUXZk9Dl4PRPjDv1S+pgLYr
G6IEV+nllh82hjda/K0mYwoHNApxdp6eI4nuKtnUbVfT8mTSIthLlhMDGeQnWv0tNF09Agg1cRog
625RzGkDuITVkmSRcXpnCUyf8fRO2VBSC7e1KP58W5p2gQLJXgpfKzPgDGqDMpZO0HmFter6SpfB
KWrvYTqkhL2YDmxhKrA8Z5yCVKn44SJ/loeq7dzWSbu2yCuHEblw0OTnZq54uN+WGKa/ZUSi1Fpc
VmT/1QDel/r9p5ZeV8pLa5tv/0a8nlA7r4w96AajD9LpSLjqmfYmT9MWPfucr3lcpNvuvyx18iiN
gJZAhmPmt+FxCNj3kO6X9T39oaRn7pfOv7WdVqDvW327HBmlctcha7OL/xvL8tx2Gy7FrJmKKqjJ
dTwmtv1SINunZzzjlV7pSQ2thb0om0oOvtCi8KadtwqMYc/oCGFZSBSTuhzREVSKPZOcXqqZsLHX
Z7crgJMsBaf4jhS0CXOBqJxGIrPzsU47ZBxBpT30CzvkS6s8xUuW0dXkEMCgmTtBBcZWR62qFtnq
LOyGEbDHBleb+rgOiR/qMLh1IO59fQxtGsSFE8QOKtHgIeLy6FzaJLDps4qKI1EHxR8DVt/bINJo
2FfqdxbRLMnO6UsjJ1/gP1I9ahwMqqhs4XcIQ5/9nzRP1Z8/Ir8ymZAwPKwWpIsK5qPLMPXzh9il
+2Y5l4YFAJ4FtKy0xcsk5nCPFE6Y8QCDN0C/7ymcESUD1jvn9qNCviFio+bM/op5FMZLcCEG+kK+
4Q2anhBddGrrfv8UM7Ed6WUuZDNc4LDAfElf0UTClMbNBJn8pkq1rlFS6CgTGvOKvoGsXy83/GJ9
Ant36FiCDSuILoeo/NZphF3PV6ttHkbge9ofNbPGO50y+kexGKS2krChlGi07hpZL4+ojUnoRoMg
QoC0W/0q552bXd00Q8tkl3Jt+mxjRwqfGNkkD6+ls+gqbQv3GTXyELTlvzbhEAk3QkrCK0TCM1TP
wC3McfzLhEon8g5O9KyHhkEAFoaaAgKquYrIbrkDh4auhMdPP+B51sfbJs3xDh+EzbPNzLRnniRW
mSB1fjJn60FXU9IHgbig+emxR+MF3xLyt9CQTHAT6wXPBXIfH+Iq9DSGRecZBFgf9oMAyqvW95DM
ZG5J5hJiBR5VSBCKmllfHVwwx04NfSQmurnqbWRrMgoPbxEfcBzEkqMU5U4r74tNfPkBovBFSzAv
HCfZ9IxRTHj4sAd2ucHw8KzbobOyEfb/Z30r7vHk92mDCSTJY9oIjIx3IdLq8vAaY1F40C0q19qj
9dorEOl0rbvVe1GcFgHBIM3xLU0r3O2RfusHpCyvVLHOfz3LuH+Aqr/+v8la399fLeG1H9ivhL/K
999PuMW5KX9mLOwMHcpa7bS6WgTHTbuxs7i38jMO23cS4Z8xLxpJJqdUOubLyYqn9r70gsnwzNHg
0pE8kXp4H8+ajEaNUplOaSrHRtmQcPhIqhHtj/J80ajrSzMzziJYb9QOn1a5YbEOljOfltYW8oJ/
OtWBmfBIQCNXOFgfBqFkCGkMUWlEBAuBaET3zZPqyKTjrLnXJ3oiVgXlhPmuyPxMJTLYmeQU2BDf
81J8pVQRBlSK1nPXCfMUGUutMNOdHkDPKkg5ncIbIWKOhm80iCh1fSkDgLJ04tcEOz3PhibasJ3C
vn/bePAB3Z+95JwSvxnitV7XkMyomgKFeP0Wqd9VDpasIw2yduIHrM843l49iuJwg+WeZMV8+PH1
K+ysjzIY/LEv0s5lkvFsDClEotGaWwsI85aR6CWagkEtK8ud/Vdf+qBYVGFr0DfrBUFzm4ed24in
LXjJJOnf/Un7JKoWXd+qfSDt6Pllb3WGYORM4JwN8h6+aDCfPurUFdMgUVnju6zgGjCIYp6/DN39
NSE+6944MJdwqedawD9kMaWRoasDt0byTsUKkyCmQt1oo2LQfQehIIPLIKgQrS821qdhT6udXxFa
UavcFF3NUWnWB3BHGHrJyRLIeY109vEgyk98dtYAH3mjhkS3oT4vExRxDvwmjel71h086zK8InnC
ZwOMjivGB+UAAnjVkDDFVmCer1Wyj7UABdCrs3dnGOyD5VEOfGU20mpmFRMTGrzV9OFhR3uU5296
5J22fTOs54LtnXpT13dTFXeALzCpjoV1ClNmNK/g46lcCJhue3VYwdbeRQLk+Ml528qFwHga+JZl
qOBNNw6/pL1MembCuQOS7PBV9EVtywBcIO9lpt6HUOd6rmNtzEWh9/uJzKzIayICC+ymjRnbjgXq
OjmY34Ym3d8IWJ5G05swVQ+iXcUelP8ESGEpfxptoMQnEN/7fHbt49NHJsF2CO8Ie1Anisf7+r4b
LqFo3rhAes+qn/Ul/EFQY+VmEkwq4e0fbaHN7/T8oWCOBTuQqtsJRhQYVx6vcL9VT935CWS+X2/D
pa4ftO6gYb8P4dyOKU+/y8sjgUpt9eQADl8Nv/mAypr6pYKtGgzQD/E0G99Zc4qMbM3g9o4FuM3/
7nexwQ3ssoFu3YSF5z2A5E7+XGte2EJ1P0JPJXRlreJaSxOT8GFm2MHHxDBJaoCB6LrH2kuVaixA
MgnKuq+S3IbW6GeAr9oQyAz9KQeMeVEJxb56k387VosbCjnKCZa2u+Gv21+zTFrAGq4uzDNYlW3U
QfbP0Ln4hIyp+IZXBpY928/M8yUXDkycwnSSQxh+oO43yQgoR99VPgnmXOnVNF8Dfz6XyRekShVS
alGn4ohiWTCKyZ6dnEVYq9daEt0gtkwZ3aU/LlL2r8Oy/V58EVpXw3rppPinS3KWlIXNXMIsIZ8V
I0vZyBk9nP63SgRRpDAVexlAJ2I/W8YqD/npUD+2K5r+bqUaXISsHoUYv2rLMiYYYQRK/jIC5iJh
h5lVc4TXaEqMZKCosuXEOeuUEsOOQHC8Jc5b0YE/fT05Va39WmDgdyuQfq1sE214UBCJx5beWTcV
rJ2Sui9krq0LV6ZCS0OxwbsI4ZtSVwuREnGtLdf7H5UhMs8KRggtmlWS3VXtj+vEqTvv3Ln1zzJU
qmMTAhWWN7TExh6aoKjCMgki6G/krVkM+qvNsDENm+xVtIgPAEjaTQV2woUdpsuNuksMcyIM2h1G
6PlFVECcX3SwqWxO6elnh/HIrj+gOi+Mi9H8UsUQuQgiv25V1M5/tuzyh2xVXQNiCJFwG0CYx1xr
pwSBW3ZtXyKbLkCUDo+DkjVmp+6x28WySbH9krYEYVj8T+XqRieEjItK/K/89JONLwJzCtTffktl
TShOkXIwPCU9i/n/JkWSv620XUkePWdMZ9WciH4MBhpOExKK03tYjTmM8YZBi5PouvmGnA78wdht
i6PxjHnU7dvgdBiECRLjW9oUNQcAtNMxfA1KXcah46nbZEp68+3kXoHq6SD/ZXU52DIaLcGU48S9
WgIwHpyLUpDs0VosEt113HknY1d7tu4tXNXgx8vdnugJZ6z5kZTSDEXhfqyCOrd+yvgCW0unFNNI
+Jt3vv3i8QM0w4ShHFCwBxjQhxuEunlCVr3kCOdsQAooViTHQB+cBzZqATlCyul0t/GEwtZAwFcz
Ftfl1BTMECtlx3PTsTq+vz8nHN+lvtN4uBh3u4LPyY3sEwZnLeuX6FF8cyZZMvbyy79qJ2D3lrFA
WGCMhJmbtYCT5wxObioJsvtRbY7GSiXM5a6ZgF9IzWIKhwpdvAWUM+KRgocyq6nkoqty5SLLCM5X
3QERZniIHFkYpXQZsEJZxws9oIeJYmgdAaDRl536C/iz+JbPiBiYXVP+RbR9Gh9uV/5CiLGm892B
0veGz0QW07MghWefh2qjKxnouXSoC9d0pNJ11RXsZmmGQJhdg1i9VFWcrCFMbAGaSTN9+QPYkJmt
RtxUKvufIAHhk00fhjYam3+OuVp6TXPL9YNNjpzf/yIRKBfN+AUKVhxV//VEZtOWXwtXgnNlNsrD
X1eLxbJSXdmZL6vcFuq/Z1UD5dvcgq0a1yuctk2EuDhriK6vw3Yw3mb680/RkqXiV/+kTO96XDZm
wh1lCQYb77IviJkYJdZjuQ3dcwRKgrxR/Gu4957XDm+UEVObYDZB7VJ+lgn2JSGiiGdsslWPKw+M
YtTItAZnB2V6CObxLtY8xwbuY/Q+eJM/JqUWbtw4B/eDOASuQLMGkL3ql0pQqmV8slH0oyLLCNCr
HwUhP9HmlUidiMNINMnF2F8zJfRcBUHwFBxIXxxTIrsrhfPcQ+lVRoL8Z7H6a93/rW24gFNm49vb
J4gv2XQeF0jvjW213QAdMJel1e4TMQVut4ozmsRi63EModCRb5UjBs/kxwQ+eJmmfCKxkKh3vnRO
QFYJ6DhVLpaXSbkuO4tLgiUgAzJ7DWrYk5gRpuwDpw7xAr86YZGLKLXJLRBNbVC31ejF1bdCV750
QwN9arK+UCuL8zZ+ljykiX4Dhh86aqXEqjh2VIKdCOjqBwN7zTIG1NUGgGAjfckxDxx3V7HGnveX
tNcg6fax1VMBfyuWeRkGEsACFC69eqBjaW9ZM4ABDDLx0rin/zJNzzDev7G+H4jh+22FMLv7MDa8
v/GCJUeAgTcgnHC8tDe5wRN743NdxOzWxeM3xXbZrD+vvEbUWX/snyEskCofg5rbuqVswEYaUt3b
h1rNU+YVY2tFGElAhzwGAUR/XLypO0x94nSX3a5s6YvjHSgZBaKPlL+lxzav9zU0sc8uqNZBZdGp
wIkyud6un1/i5isUC7X4LfPNB6v6mZ9lHfcOmOhtfck2mwSalEerQ+EfWs8rrn+V8hUg2/r0KtV5
EVbJf/phs9cuL7fV+AY/ArFxluA5JF4I7HSflqKbdagB00+OMvzgIEjjMPnP30LyylYVnYCoGxtk
sJW9sSq2Kfy9pRr/anRRZdOhaYkMuSynYr6b2ykttdC+vdpZtPoyCs9gBJeHPsKP18vkc0TZsaKe
jWcnsCjSDgA2pUV1N5NLhSH6sTw7kJ8KyrDuBRkrC7RXVTJ9yVnqIPaL3JN76nDeruCPtxkCz5GX
Vtvw+3rsFU+8fQsiRvTAWEQi3GwX/rSmDjhXA7ds3uYkJAq6Y04IWCYfdzsYPZ6oK5nFvjQ6dI9L
i9mGIHZ66qAHhzY81S+4jbAjka/WilKKBxpuUxBPkcqsFkD6etjBHrdyCX9egVlcAullIm+sQ/0h
BZJRjXJmp3iAC/2JgWn5k6TNYbEDx7BYLZbcIMyLxd8iojR/ugeKCuu8LxPrEkdNgptUv/H29CY9
8o95EUrKJw+dUMLVtPrDYEFCuHA4wU63Qm1qTsZdGxw/43k7DgYe5Wl7TPw+Hqm+yy5U2vGdjeEx
nd4kOvr0r0kUIi2V4J3jVu9tyURRrBB7j6loSEplFGcb+4GBLK7D6X9Ai36/acmXurZ4+qIXxI4o
98PBVBvsmCaH1ngqlYmu9ibjfzTlbsa2b1jw0MilXqFd3bevQdRwUISIfGfdiXZtPQs3MMuEvAlI
vyPhkBf/kcNkhJ91pWW7Ddi0UhdfYaq8agT8X1zlRx4Iku+DWdnqaNYuGoisNANzoGOp2V3dY1jE
0zfs36r/Qi7c+d9je+RAEmC7jH55Wd4N0d1EsseVcn7H7jnIAVHjf6/9bI4JGTxK14HuOtL+mxy7
9CO+QOOM2l5SoNU+XbU7kdmX3XhRywBuBl64i68HXXrdsYZy4c+RqxKW/R4akf7OvIOHkDvJVima
S99YTfvWJFOe0OIV6Fu5vdcT2nfV528Sg+Y3xHbyn1cQSo/OSFmafen/SKq+T5RmAGVn1TnMfQ4a
dkGCgumI/nowHuStr7T8Tk777sLXYb47TMZe2Vbz6LFAvVgSnINGbyiPNGd2wmsHP7raYVgKHhKm
nfIzHRJl45TpYKEyi5+3RvRwpYstjBaDAlrUKwpuyUIsaLHhf+9Zpwr8ixC1/dy7JOfBs+7XnVT7
44yb+pcijmKsPwEvScuGNdrcJQAYfwgVaJf6l/nDhEfVicHwWkqnSAKoPYs2mHkFZB2v45cXSawQ
iU2k+aK8MMEjJds70YH4f4h0MbI0To5DGdXmKYsqQkhf5mO4R93Ms1m0xKJXIpYrv331bbKUpy00
juM3SbwsUgaOWJwKfrA40hGTaKDk9BCGVs+pwxCt9yfY2FvxLvrxek2V3fthkyY1ujbh9rRtLbH6
hK+uF++ZzVEO/fU1gFQSvUZsFqSboeo0kwO9FxEvUxQrhDolaQgBVAKgxhSdqEz5WcC6ls0SdSew
fPqKdSkk6QF0xFUCjDqwblrDkXlq+A51zuEOiifLW/6sxIH8PbQ0dEgVJ1iHPAbGu4uFwf3k4MFh
cjAH8HVknxzTpTGZnl9cif+ukD2HVcKNkigflVhwPH4vyRJJpT7BUDHAy38vC1ME4woIJosYRq9Q
m1yHcTDAmtwZimRHxe9hk8RkneEq8G+0oMG/6pNhP/sD+aEbBfKu4vIkYSDjVM+HI3U92Hwwc2gy
XiBQ0DB6WAJxbTM8Xc/FRfm3N2tnTIUhfDQ0UoycROMS0BRqGioBeELnwxDXmofZlZQLKFdWX2yh
StaM5L/No3igtvmGHeKd/Zw6awKnInFsjvum/FYhgmLqpme1bZXH/FQYxEzl/UGAceqRUPSDvkGq
ADEymS7IM5xv0f9jqjHmHyuaLE2cft8nR9sWiTi88G8GQSy9t0hTZqE9v24HSE0UiwB/1e9rRTO+
oK4/i1Z4WwEmUN3goJ0BY8+CrCfIw7Elkp4BYiqxP5pCyHoJfxj5dx94o16astYS4kIC8XWIeB/H
AuFqOxx8dVLIqPUsjarNxd4g09YsNmkRNFVRd6r65HLrPRuxlVEU1QtWy6eiJHg62ksX7dcWVa+O
dw6KB+kumWBe8ZRHzFvi8i9q72Zw4gaefuLIfVreI8aABKWERNwPKhB/xrO3ARukoKymcSgllrpU
AJTX3w4w6erSNbXErh9RRjmwSaCf5T07Nt87CxVuvpmNWMu7HG+Shp4LYwa77KavUtGe//APvej8
/spI4fwVZPUKzxSMresMB0u3DCHba7Z0NpaYqXK7HeQB8ST8AbStbSt3eZpBy9k47hNWVtm/UofB
ufgxNdEoXBmuK1duBns5I4q7Fi4X+7GBhtVe6v5t50hc6aAsZ/6cb8js3kv3mxez/FxQn/173Loc
nrlKRJ0mfpX5rkcFQImjVx0Flc1EL3MMDcfadDYDZ9b/5HL52X+aifwFsKJBCxV3tXJSxbSXOYYw
HsYhDJXgESAwJdecMcOGC8/qmRdm+Wy36hyXLQKy1I/WFq7gTeGRc5QCQ6Zbh4KNuWnwz8fF9LJJ
k0l+9LSS+wF+z77GFzhM8wW69cH0lzA5NNIBrGvZkgud2M8pap9nXF0cQuGgVKgCUoB9/GEFnAR/
o+wLtI0TS0HbKldZt/jL9mBmBv9B0nTpexuJdlexQhxZwkn0X/Uf0agcy1tpJr5DFhlw9kVZ++v6
IADqzsxXgCLmhvm0y999oRd3hVYAm6sfcIadYzeVeYMazoX381yJXix9tYJ+vhbagHwP7FN13++T
Y7cW4Kph8pMGTol9SPFaHwAt8w0YPNphPAGuQWvdLf6mpXsZsWk0g/XktVMdsKXILuBCbPdfG3rh
3e8U001SanaH3mLOW/ieoC2uoZgDIKsm9seQgJWaHYKzmA0xlHOx0w4/hkWA14JO6HVuTan8lARn
oW8joOWsxw4X09kMoAK+c+zJbFlahFm70ldytb5e05q0jeazU8iWk9Z4xt+FrpXI/ADKKIpEEA77
EEvRsE6XfVn51F/PwfuFB1UF7quTFQBGqj6yL+q90EG/LA6095CDwVZ91K4uNSbhr8KEURXB+20w
VVp8OhFlOBQZjRQNcpVRHddgzX0JiqIrnzte1J7pk5GE/v3sOyGisrF6bIm1WVjFweMNkxVftaDp
GVL12Qf7ImB2d3N6WWa5LV/Qb0f95UWNJuwwQg/PoAOTtN078LQC3SouNf7H4unFrhJROr+qauzQ
+Qr8IX8VTBwK/lxKXWOIRABN/+6724blbZrwyyHUxBNWrnU9g91UgCinREeebMHJpbqMenI0+8iO
ImyaJe4krYu9ke1un+TyaxKrwOUSplTICCSlzpppIaZnYUdKX0TOuVND6E2x2x8pk48V2vQmugwg
hny31wBVjyWFBO8zz17Tb4P4Q6s0e1rNRk0dEDs7QtEBHng8r0JZFM7jcUcJc6XRSyrlU2h5mAQg
W6cTmMnQuurjTjmkUoFqI/M/EF/Oa4G3oroYTBwECp7U3a9HeXJFRuJIympPhu6eVN9Qy4ZDXxvC
gzqvxZGmyzQjXW2H3yrP2wsJXAHV1Ad/qCzvjd5NzKCJRaY/FS3uhjEF8PjFPL5Zj6Zn4CbG1gjw
zsXh9xITZvF0jsUEk7vsZ2gCXqAoYgJ7kQtZcL3+zWrbQ6i4Fh20D+LFeNPYPj/8a2ozGIuEXIqV
kySRcoLFYfudYqYkuijRu0CL4zPC908Q7DRDEhPwnx88528KADXUp5RIep47v+Y9SrSHQaYHWakB
aFwmuzFUQZzkUr18xX1fIoVzmm2SE8ZlVZGyPMdfvLXAwy2Ir9A4sTB3TRXky7Dwn/0L8aRJnXDG
Tr2eIOuHJR8sAIVGmHXAwmpRhXtIcnRJTVzXZeTl3V3vSKyfrn768I4KxDCetqZ9AYmzIJYsFzRl
espznchdJN2T8yZN+4B/wIr5qRfIQGUaZcMyxcaxKFUYWks+GZ+jEYmTX0sBEuZcZ8Bzyx4ydAsm
wr88G4he37Rckd3Xv7T8iSDnkUA+Cz3kOfLhjaiLwzE8T5+LBoLt+HSyKlOZXUSQXfq+FCcaqDlE
MOkJYC+SeqFozgpf6KsScheBc6Ojt8cHvJJqIdIS4p1nMmh9XM+DbmXzlDyzoIFVrp5TnwZUllWq
izHcMwtzoW/V3oWcffFrLTrqwKrsgCrgTKzQDRa14veLCbkKE3GxbeLQlRGi9vKhHEaCEd/VO3Y+
VVckRqenmtuHsPNpg6DKxfFBROZ9eslT6z/d/+f4ZDWU023dty15uMPlnwcW5WHe1aAEmUWYJYkS
jqsD5ZVyBDy2H2Bi7PZWpytj/4TbxkJWiFNgkeZUF9HdVCFGF5RkA97lIc6xvxgSKjn2m7veQ+ff
vPM5ybhjejKk58IQpL1fSJQT3MXg/pnUlZMxVh3cRJlUvHhiC4mcohVEts8K7ZV9KkdGDBduhLyL
4E4vhLAEpS+7C7vaDjc67ARxZWTjIXwR5GbfJ84JZVSmk6Vr2DS7wNcI1ZsiiwPSGExdGjw2v1gp
o1B82HsYY5jXYHUWnM1AEzhhDP4fqjXA45aiER450Ug3+Xh9siHWXx/LRXDq0n+2UmaQv9znZbF9
ohHWYxrdC3jZh5IZg7J5WTk0fRVHrHvSi9r/Ex1SyM2iM23qVVqzfENdh7X/dtnjR2Rv9BCOLAN+
+vUA3YIwZTaEZSGUSWxHpEL26BP4H84hihQVqLOw1hnKz1Z81sxfUEYkvFntJynZiw6SjIGy1b5S
tJFMc7csHMKh/+63TH9Txm55ddWWnLQhfjjhF2WYzS8IoFirrpsUrlbNLPWmtS09hXp219YXqpBG
WYjUfQn9+B81jAATggCUmBf81jaFM4bLb0uYdMOyglbUeu4a5f9bs730RzJ2divyHaHm6VU9io/S
T+/0tPC4FmoJM2knBFbKpUAxM4vepVDT/aVDekVVBDhGOK6aC8oBsOPnLAY4ieQEMS/HqNu2ktCS
+Gfp5CHMIvK9l5ilBpi+zGw3HAFM9UIxaj+XlAQAMKsMpAKLzRPGGkDRVOtHIv/uhvDizOTqg8Oz
wJ0NpNoEaUMgh/OeiX2i16/Fe7Mr10wAYWQrXSwi9kpZ+myTqJcJCZptuFziJjVyglu5n0CTM+ma
9Cl0Kos6UAKbcVZ7cUNDL7uQbe+R3+ZdvMVIFhQJ832Mn3chHivIfRtYBZs7zEYgzk0uUwMeqAcd
wWtMyCbt8/uZFEe9gGwl9NuVgaBqK36Ac+XtdlABj7UT9QNGK7iTwc/mgDz6HS4oiVQscXxY22U5
vTvcQuiqTfDUwcWtL40/YA3/sdUNmvxxm46T8/WTh5luNbzOB8dZdk8w7dbGLGtIWDuACjsTjVN0
ZULY/vwRWUePr23ejMvgOF+p45mQkfICjIzm1vVyeiDoHnppAwpgWk4ESX4aR1QGoudpJ0rPPsYn
uI92MGj390R9AZKRH/C/Y7r4TD19I/0xamgq+2YZviSG8nSe0aVBAsWdln3vQG+8vZLkDyoKklup
9S/stwzMyCRxn2rtM6GzOCImbEQiYxFn6gzvdvKrSoJXFlbnwh5cCSZQ4a7Rm5qxD63l2uxFLO5k
7yw4VcTbh3sCgOAbhlnJGC0csaWWCWF+lv54R4q+T0SI0yJY3+97i8ukxmW19h3O6A1GABrhwqoa
EeyHi6NW6+spMsSoIAneQreQVfTHn1U+lRDdyWFIyp4dCCgRKT4WPa/SjjfjBBZMc3yxbjW0BB67
32tXzbrw/dSL9rQppC16CvGAziS4LQRezXMsKx3Pz7b2IGW7OxyirJ+j/ZdTbAl1lHSxtqrY1mOC
0QLoKsTkZbRWbKzgUFopQpemalDlTxaC0x1Z+jOg56+gsfoldZ0j167MPta5bq+/qocS3nx1O2jy
etfJECb1ZZluSA5U2e1D74tiBUFz8ST95JUlBX8Tkc9EqvZ0K3Ix7C1pSzLXdxZDh0UXexe4+Tnw
whRQ/HejKQ2/ytytcuodUrdqKOxZk4GH7dHLmnZSa2MPgnfUPOwYhoT0thPMGPP4QFWRzms1uRTv
GkbB7E0likPj4iUYRaygrmfO5z8SgAtGIgyfh4dL9eol0fY6dPYhmf8KBe2SK6wnSFvZc8iEYuj5
DEjHufG/oQP5zKJy/YN4XrmFbEzgbIwudoM5WFUsa+GfcJCmxuzmS76rxUQVNeGUJO1jYiwAf5X1
XUYaSYJRq3uJs7fxlBSsaQlvTbVNSqkG/iNAatrDDSCEYge8GNykJTeXWRjfd7OmJWDlV1QrRYee
ouuedyIcfE6SA9CqvlPwu4EBX2KrJYUtLfSttvh0F0ae4GxB0RFwytnphUPw8H0OpoqC61PUCL1X
5Z1iz3tk6Y94pAqw52t2ABcqPG037lmqX6UWKW+WTR5fF7T+rxZQVD+BBh2ZV2RU2DL1OYr9wosz
hDboFbHagQtKQv9Wl1lWHlSmWzNo4Xt46CKFI7dwf65ruPE10vuXh6aV/TtGvr9ArzgFv8AG8VEV
oabjvzqPXHH4pOQXMLbbUoOGsmeqT6wBLl6inSXyu/LjURaO7z1gQkrNazhOgq2XKNxN7NWNhfy3
SKTY6AMMhIt/GoJxD1u6b/bLgt61vbRKX7YKygj64oJz2q0cL7S+/UULvDtUye7H6tkOLk2U3Y6D
+whB+Pjc6eud4ZqQZxCY8P0F71sw3s8r1mPBHDSV/1PembLGfuV469/i59Fdb5xhjl77OuU5N/uD
GdahoKoJrY9UrHY711gbEAnYFAd/jm2H7OLbiIaxKbDW9rPtQcnvegapLkoXIy/35NiReJYPi+Bc
3WGgn1DxgHdJdbv35kckZtjhAvsZWOP/mQAeLcUvIYW/N/ugi+g0eCH53MFTeQizlv2q2Z8XSYnQ
nMe5p5cX2OR/TDylvJTk6KwaJ1RFNYZlrPh5SRfxxiVEUF2H4cq/7duEn1OJRO5RnTUiOa/E9N1C
LQG23kY2G50q4BGDBTvc76Tb+HQQWj5PKq3TPdX2ByFeK1i9RJULC0FfXGCCnggiJJXQ7rZxL9C9
SuhCUNURff/9kRbMviJbZ4Jg/S4OhpANwg/CA7M04NYiOmk8X5OiyZJ+Q6h4BW1DSbzTAmjK1qPl
FukDcYhZS0w8AMwyEyRKGCE8Ds16CDoUTuMhxugIJ4tJOWzT2BdN/5k7ZrL+eejt2nUIPC/ivSVg
n8BQo3t8q4J3QpxV+XLuOWEzdAdOkHkieEft63U+8j1EtUHpcsSyw6aPNbQ262OSKvCtyT/cMFBl
rEOtpfR+CzpYamQwTw/faQHi+gV9JzJnmt54yJTRotVAsiEaofvSrmnGf5GYQEA4zS7JaJtX7yA7
QVvJKFgt+HbDv4ShIaFiHqSjBCMd8dhO8368RPnHBYjYNfmwPPv55XT+U6YZeWDTEY/FO8/vpLMy
2QwilJKJs4movp5hDc4GUxTC5F7EyFboDPDguGseS/9PAkIRIqM0mSuNJxFs6y1nbm5GRX5Itcf3
/DcG/8DO8zWEDaJK/r3Rm+tdLu2DlBv2Cvj2fSsiI8oXj85ofqHDe7QcbAo+lPtyTJ4zXeLZdkC0
klHTig+wKIj2+cZ/VGf7/Q7HtEIL13vVcbdZ+SckR4Mev/z1fn3hXR1YbTk/5OSAllLkjVYnOymA
hoYQVQGuiR3dFvuxz/pjlSe5BqMDSOdRWRjg4qYuqnK+6AwHkqs+szf3bmPWYkwApgBMOyxGkwzV
G91nWPtQnnWUwDTyrhZmBIil/dd++VheVt5OAqO0EKEF28xXXKEVGQTDZHSN7kSKi45He4pncc0W
YCiF52ylii6COjGxHIrdNSKUG5/MJu2510ocAQUumacEkR6Xm7vZ6hrf5KmL0lJcq1VZObuI6Bpl
isqw2+BMQQDWQnvuNf2a+rmeJjOmawRmuQBV3WcdVKylN9hXgSgrozto/guSuvbb+t0Z36dzDjAU
fOprVFOrIEGyq5fl7e56EdjKgAQUBI9x9Yt7GT9Od3HV4z5kyx7Aghd89COHD8WEdr6L60m6hm8J
TcOEqLHmlAvWpg/htyNNZh9NMzxZYsrVhQtqoe0q/A83xv8HvXNv67db8RFd14El9RO1yBz3i4ot
s+Yo0T9T1tLQhZqv/QoUBnBx7zL14HqTAnM2Gtn9bJgtAwOlKgEpYwi7OL82aK9UihDKwsniTCaX
Rs4XdChNsD26Pj/Gw5s8tQQRudhQp4ZzYuoE/5N6IRQqf+RdXEnT4c/S+FXDcyTaEt/TUdWcnqrP
+CXn6cBxGPJ/yVnOPkiGawQHXbUCDKovZHWeTjFnm4jrbET/UrNKVbsRf/ofiRDr5tNWECsQPc4X
Qrh/Kzsuxh+ImefxQNoLX3tqX1PNzVcUZJzIqoDFv/3piQlWvpijZUxQuZo2sE0CElUqtKCo3k9N
TegG0X8yWBM30v7QtdETzIoWzbSyQgEY1t1EM5KKWv2LQrnPietJ9LFK4jfztjkn18Yd+fMEF/OZ
sgRyFX9PYzVdqZUAfaC40atq00e6o6J/n0gU7o0BmnIDIrvxDjZQzAsOiQsm9f/lTC9bRIMSN7/H
Gs04iqgSw9fWwgQLR48oezNotwrWt+RncijdJE/h8sZ2CQvzQLRpdw9KZVuUwsdgkCS9DDrXF4qU
uLXi9qhWn/kEaIEmZada0Kru2KBtcFAyUjMc2ueMd5eeBbWVpNl4nTwW6Rrv04VoR+osHAt0L3tH
dAt0J4GHyAvpXAel9He5cgBeHrtT3wJvU1OOiuB4FagaD1rP7tYiPsVi5xaYKtwMURw7CfhD9W0A
S7Dc5mh2s8stqDozaQUp2rERxvnmN9dmrd5A3WTcKrpUq2wntET0mKau95WfJY6fqJHcEaI0tvWT
rTPdhqy7byNtNuMaRY1ytbU8jCEBSvwzqFpeRR6GSiHTkmMw0Q3+o7DmvfBzvDO63decidm9a5SA
NkBt4As5c6LdOCIBjQFitEITaNvaGNPFZyXb092obnm+5fMVRhb9cqj2srsl2tJ0BRPVseF8Rq/I
yQWf7cxBI/6DEqZHn2yeXIF8EbjachyLQFYLsCVrMSbm4GxYxeBx3wyzMez6H5tZrhqeFhPip9k2
zSHazrHayBiUZ3PtlGow9hdVh+cDktVevDwl3SxFr0zjB1dGtwcU9hePPk7WC1k6zxs+s1t8XlVn
N5g4AYBngnckz6l3AUIaE8NDpwjZT9QIB5WkxbY0XZFngMJqbOzG3S5zUduh/Aj4R3nZVlwohc0+
UXnOGojMP12JrXf3AuYURucQBGh5EYbY1GJg29brpfSWqEYpFDEOb1NxmaJzqr940HKBQmnHDhM3
rql9s5JJIyPS91qCp2nhP5AOGXNmus/OmlsBfpu2l4ChpoZXcJCX/0J3sUIEKtIrZpiK52OZjBZC
CVR9wYJ8IZLSH0ZfV5oiEYq0Sno3ibiGS6XhCM2Gn5DqhOiMdsnYPv4UY9EuJuuLnlkXI49u5s1I
ukQXtRMVVr2FF4i8OkLUlAGb3RgQcdt0hRUpVWw3ylv8fZtociQOP24OcQgFhuMtT6kIgsRtW7NY
scNWgmwciorn/ht6CFCRC8sCm7pzDcldKxp3w9plKSIsMyqL5dEDLqz80ND1By3UQQkH0nLldFj3
ni1DdfG9H/1h8kYYT7PQnY01SHJjs79/xgbN+xJ+MZm61t8M/uZ/MZrwGhQqnAT9Iic6vBOAzSaW
j4mjnEHELQIQeAhOeOYKYm8WSGnlAQOqjw7kSPv8QPDiajJmj2OrDObR4r5RtvJtiTaORr4YCJtC
aDToFASe/b+Q20olmaGPfm5Ri9vuisPRSlFrXlblK4SGwCfy1Aij+BwpyNOwRL6/TPhv8X3KRR2G
SFWDewH6eB+LZZM27a4uPUV8/BC0Dlto3wRNIqe/f/KhIwSlv5Wqi40MPFICOoUV5vIwtxuMiMxa
xofxhCkcVJLFOhSQZ+enazCULgfbxrjL9yzK54AOb+hHPlZbgUCz7ObYzLxWbczh1CZ72X+xNO/d
PC0UfE26HEUUWr/L5sZ5aifxgQuMSE9G+vLEj9nyB3UMaVYd3hIvJRKux8xrvHtx3oc9u5/V5XU8
ED/6XFZSwtTLR7zk55sh8SX3TLUkovRvbNpVqGbVOXCWJ0UWmCaQWvlfNE++t6JEB4BLXwpAwEr2
E8DNJAfNMAJZYeq2fZ8J86bbYlJx4M5sC3yxLSRfKo5hVaq0Vq9UMmbXOTFTHEdsZ4pUd4LtO5Hf
6EBjfqu/U/1bQmQR7tbgS1QjoQpQeUwMB9RaUzzbXWecwYYCzonHukEJQjJHnznhhU63XEbu4OU8
AJtPqBNbiNuS/3AkLH2YWfPmU5KQ6KfS99ofXSdqWIJ2/bHFs2Nto5XJwA73qgjSJzNshfzQW8Wn
NAB9qJzsY9u+K3teq1ns2Dlbs14HXCjMmiGZOixFm/k29P0qwI29w25Ue0f1GlsDyJwwUFfVbQXG
p95SpaUNkZST/6gs22W2NseWBy/MkQgtmwCEkLJEQsNMurFqpKW2S8Q8G5X8ywUWvHd4z9vE8Smk
9xvTeBIsg5OVYWjBXuU1tGuQED+kk0TfeBC7al15M8qcOrt8TBjV3JwdoIhp7+RcNPJFS8cZPPBH
cMPSxYlHGSDKL9ws7SM3IQze3yq8zwIDOEvKgD2yPGNKEuHZ+IgMoyJdiwDHGLH0q9qZeTtNgSha
a8yxW9OfXAbnvfJpHWFo4ntFCrtbypgQh7roniIk/3PqHGvVbIyDxeSsZ8JlByyAhDDboLeKJp1i
wn6XvrGGL6LVoqghyYmXDpZz9jE3w66IOst2DlTLpUqOih/v50oQK4Qu579Oio+22WEpLecUv90d
GRcdESYJiNtsjKkikTaDTCqmkLpPr1xcqyU0NrF3T9wiSXzFnss7heM7tbPH/ThaO0y6jwkzz610
hrfBEFqjNzh8Qli03rXzL6/zO1QkTwxhtCMKaGUszhAevPjWYAWGQiysO/T1FZx/h0PAIccab95C
qD95mpFKktP4SZm25sAO/04ETIUOsQbdYRSIyqFosQQkFjNwe7oGZ9hMF0gM0WNzp+OmvUmPAcs9
q0kqrvHimjjKGE4tTM2nNRemwXqVmplj4P7SSra0CVuOHkLUmWEYlblfI5/Hby+Dl1gNeRYeUP0p
lZhb0XQezlDQov7aLUAcHedMe/Bbkp9DmNFhiP5TsIDSv4A+KoQJp+LwfSO3lH4Qs88nLmpHTKSg
upDoeFI3vdpYvySNTcpE5AAdnb/vUct+TQHKQFbae9OvnyxTrO5lYnLT/S+vPCtN7I+VybmUTJDq
Ohi9CCNkoIvRJVhU1WSVtvf0xWpQ2vDMVne3w46pAy742aIGX9jYRq+6JQXHv2GMxU7DctxTYmBr
jdZaI8tGhvz5IANyMUp+rIXIgqMBYaeK3t/f55mU0vRd21IAsg2u1evZv0zV/VqBfhresyh6brbD
uAI6uosP/Uw36UMBRFH9jisTXNzImScaKhf0r49U131YYob54XgirAQBrMULh0wydfWEqhQKPYZ3
tI6IqJLABLkh12/HWd6wdpk92rwTdloJ3DxQmrH0GRmGbswvgyxrlfsN1ZmFcb/bt1lABSEn5ku8
/5DDb1U2vujAs7gJcpjc+WqelfOx/E0bk9GbuAXcp58lUr6TYsTCq3WUt/I+pD+bmqGcJ45b0iL+
B42lrwaM8ryr64jU9vv7Oay3QUnlGbpGAWjsVBzZ+RdP6MSmOAEEhK5byQBdpZSyxXlSKg0aQoVB
a9LtViIp+S964yBgXi8rdCAvWfEPBEjKuGIsdOnXBH76+OhC8M5VgVecbYqMJrgmczYkeAfhrUpG
nZj1E+AiMjvsjNe8hmclV4GgSuGq2hpbK3CXs6wt9t5/yd2rUQ23o1qyoSSFcqycJA8op62HHNn9
TOfDQvUhr420HTCQ8p+1lfMmXKkGlpXjI/eY6sQxDieEiCNfij4c6DxHBQI+lZiWMU0WEWNUbjsv
qK7/8Tc6s6dz8MGf6+pavq20qWaIPUyQtU+W20QJKpJR3sLXef8Gvr1wIZScVJaP5kuSIxqlL1B9
FfbeMZHvBywirqagKLzmn73GwbcdWj19C+kHZNcrcbq/cBXVWXoiC/vSAxsK0SKI4izWMn7uMjbN
pHu9SyXWrA4maBqGB1qeCzFStGIbAijb7thWie2n97mpSMAwXmBJ03Xg133PlKy5a71ShKP/aGJJ
i1rdR/qdcXtZYHShibXqRTPmcGUJOW9SeJNpTNoSNIM47i76+mCn2vasSSFvuxrsWiC3nT4DKJxE
EYPNYQCnXApVYBmf9x+00Q0uw9UE8t4yDyAEv9D/txQeJJIpil626i0IQRBeFniTnvsxdQLPOVO6
rok7shZdHtOgCkUBwdhIaSov7O4MA6yhaZqiK5QHgUcpXU4NZOUGjWJxko3gWuAh3958FMErNtCo
Q3iHAtHbmSUZaglCZJbwIKxT/RpoU0wHz2ydkPSHttBSD/RYBkZ1guCAIhLqiZ0GyETwVYl4hSmW
NDDbxV7Vnb5NnEyrVO3M30WltrOVGfaPDoSxaPhq8yGP101aywDbqu08iZnrEtosKFEmFVXix4H7
WHz7o04+JscudxpHZiGGT6sASlGZMfPgTlmAI6v3PAN/LhFZUxxDMlsyamxWve/V0pT5Qi3P5kQl
FZqoWmB3ZbQ0Fhxo7DGh/Y5xKQBRRa1v7PXLb2cWOy+Bugbsu41KE8bf1bVWXpUotFMW5Tpexc4Q
OLaze+hKwwwaQLynCQ948n8/3fybK+RmWuE/ls/Hbz+Wa3c08p2j0POsj5wQD5zCXli7WS9E3BVT
+cA7KHF7Idh+xtEiPqCoj3ymEPI2C8kdRhfkx0WaDqZlaKDmZ4iBl9kV6vUq/TXACiC6gF71uHE/
bxy0B/uOSrTrWucqCmHiSTC7NPr7gSBdLcgA1mlwSKkqAokIPeSor7UJXQmzm7SVzeyk+UvNfazg
6XsieFb9Q1Nc2qKv3Boc/6kASs8xO/yCfU+fkT3/SDTVRDPNRCRr/KrsIPMcooTJA9fLjMoPYkYO
OIlkzJFZEjmPiKFRh3+H4CQVVxFo1jETs1ZlmyaK4OcuUH+cGltqT4hXz3G8YT6qe8D9bgSNxYYT
lYfzzhB/LjBpNEay6Zwv95mUErex6sFhIv/M/S/DQayLRFcPCNwwb8OH9n6CiHCgxSbzNrlaxZ1A
7+p83fxfYGKweh6S2qw3eZTmmfdgZEMj/8puqLttXlHaNwjhO1W5VGO07htHz1WHEPikhfuP850X
IfJgiejciDpiI0uuVgQnVaOgJlTz0I3mPhJFSTGRwsc2QxVcK4DZdfzbb/5oPNTUl7244yHJuwHp
a1bXdNrSsyJOjGU6pQBWG1EORbQMlJSU5Y5WkhuaTq0wBCNQpvrU43u8UaoCBSk/7C86FjcpBsDj
iqAx0FdtpvNu8ued55/YjFyRyNwU56KxMBGz18s27wpYq3IyDLpv5Y4pfoRkRFESMMxC8Xu7LS5O
rQ0s5kga1LXFAmRZvUjwCEXI6WlSBKS4lyJW3d0Q42vxI/OcGe+rCLpC9XjdNun8XgMvqj/QIMKt
qcGYjVKkSlJ5lJsPukTd3B3J6K2LMU9Qd0Y3c8ZtWjzKXulYtv8U6P4nN9PaWonS3RkSmiZ5VHxr
LdVyMiU/f8OA4es7eMR7KJKiCZ1WuzHffnnwycvdkmJQnBOYrV+JD4XHO0nv4OQ2kP/T5fOOOUHg
gzY1WcXYO1MqRRJuOytCdMQ8u2lidt7YDeBI4RWbEs6VxUy2owF0EfZSsvQofCqqHyqzzXkK4guZ
uXeFWvAyEgn8j/s/C8vxQG+8ytRwr4W5m47f8fIpFVCsHX3YCcAhHYNTN/47gThLw+O3brE+VEAc
S7thG0sdYcmT9jNzdrefB/ioyTU6g7vI5VX+UVwDVJpQWDir6iAe7Dk95PcvfOhec7K87xcy0ATQ
QuaB9RANij97zTUaY2Zzw1Z04A3ScVO8vp55j/T83yc7LqCOgK5YUIKSMsPRxtFBlTn1wZs9TH/8
9zmpMzgsIlcWzduUI7ML87dUSSPDzxGkAVn3eacedOZ3PGInZknpuiTGst+mIkcwOdUAdDxQIgB5
ltd3mZnKJW7YdqBDrfGXMh0IucE+zm3k2al2MtoRhyVxw96EVcgt+ug/PIi6ns8b6Ymg2LgTLTvI
r6RZLUu/RMQPKmiQrBO41pXtRUb4r8iOE7XZaDTl3+D9BCs1/UZwNALz7eJIzi39ncSx0bDTbhi1
4jAlpJmIsvlkulenYSU9Ei/d8YV78ymYfd843Q6chudvyBzVhVcxjwA/syCkAWoAS9FQc9rDbkCV
4tV/c4aVzivpPh3sB5OJ/XLqmzQy3bOkbHIqSWsOqgp3sc0XNlNuXqkb6HGHthPxo6jwuTIBv4Ck
rSuWdx1ZUzsv23f9EGI3duGhTlAsiuZULQU9EiJJRrL0tdxfAL5eH/UZipqCXAd1GeDVRd8Zcy78
GY8gZ5/14FDk/2eWrDvhBwXRs2wmW5WQJ8nqrcrmKeNyuVnVeiaXJ+mk18R6tcKdQTkG/rOJezZQ
ZzPu4NQnkYXA/8VXt06iToJSYMLjxYtlZF/DXZDDfQDiFxsdyW9rvfB7JTJ3YPy54zTZsNYXm3Hm
UOapptKeSXPa774vxUwbPRoXuA1jrDVBLgu+MErf78GjbGyXa26Zfd3pxd1yLXJWQbjO6/jtFbs0
dUFRPcnYZ8jtf0aDNTZ33pulux2Dl1zldKhf22ZZszeejW3c9y3KIMJGUx62vMipxJBzWEfuS65L
avSy4pjwupSdv1qFa8k0xvkpd2YjRShl5CBv8xtlVLBJd4biF81WxmKfoHEIzAqnBa3pWIaz9ZnJ
2OhvHkeBWtjZG1gXDv5zCRUTZbBgl5ZQl/ikyrnu/v1omHVe53hrYWwEQem9ilqBSfBWNIvg/0oj
SrC8xv7GsR/J4ekZMbZ4BeE8NToal6xEH2O0/NKmnpuZ06d4e24QoNNJhltH3tMW23+V4FOrQRrR
0bW4M7LojZWF3JOV6YZbOD78UJgHeAmkJYMPY8GfuOh254YpVmujcs2xAqBVfktTeVin4Z93VtTP
SmXQHt/7j+qJx/7IT7B44mr7tfVxpwe8cCu8sxDMTnSeMFy9tv4n+T8ckTJ2qSP5+YRRymrlUfvi
dfxvnHPjENlHlPAmjwtcisyzxTzc2T5Lj6m4v6ppWQj08QUQ8xVy2ezLsbAtk2VVJEDRhtkCnUp4
+lJJKko2lS8EfjkHaQlMguCsuznnZ9k/b3l3v1llZvkq3JZRzKV/LsgETpDRqArKkUwdKNzys+H5
WroolVNRCZ0/ejscWgwNwYEIWMUzPNjxpRwDwIs2ZVx6xZpN3LR7lgv7uJ5Y7rbBhO1a6e5pGy7N
mM7okZYBKZ8tywrhTnA1oSJUhybpGuwFgStgSjgZhOwdmw/FJP9o1VIChQhkipSHddekPZs3RkRj
M7s5HmOVHwCikpADJ3TZdiBzMOO1kCwKp8a9PPcEYKV79aidO2nY7fRmRqtF0iBD4TC/DNIXY++B
IWuRKaZ1csZ25JZuaOjMLxA+CzErS6NM5AWIn1BJE7NiaRs9ReIxikKcpDtv2bvYAnb5kSybYW0g
ZkemdXQkWdL9UETn/NinjFIUaDehDdCorucHkgD6HhFekLR+evOlUhIfbIEHoWxKk2DnOvRa8fWy
7y4l9ZMasfhVjit7WAy22f5/tFXgblwNb2TW4CnRlcPrxQKdebHqgf07/f/f2K0kFA/+1A9hv75Q
iSdiU3etqXwieEDWfPIH1y7P73DDHlUXKXIXyqtP9YdloIP1V/lSsma7e9wXpjsR2vCe8s0/e4lw
lwKNUhfmarZE8DVwWOdHUfigNwRKBiv1Lpyhn2BV9Ia0ABjg1OQ/EKKtvzmozDmE4+T1gIFMx4Nu
EK1wEGKi0eaIfy+9uLJ/VcR7I77NhJ/3HjSdprHVysrXwT309ALvoeA+NsEeY0ANrRDLrvvhPO8Y
cWELusf2752Ufsrr9OCf3DnYWbN0cSccmAsg5PaCndyIuQ6xGupUSZdQF2w0yl8+O4hNjba/M0ou
cbavhhfkwujap4eRpi2I8xjX3NCHj7If+zZAZs/WQUWhuyH4ib+N7d4MHvCdc4BuIZ+tH7N0J1As
MIAZqiOf8W+MDpp9EnKW3Q2B5fJnYCX0cCwZ4sMfbnHPek0bfS1azS6PFQM+oX/x/j8pmeCRNSNV
hkwW5+cGqq7/dbImH5WqqgT/iHWUil0QZd1vY/LYQ3ENZIa4e6idbHHhkeDayhVXKxd7IwpRP0Dn
4itwYBFANtqV3UKfCTCXuP+tSWHFXv3l50o/7JTqC7aMNi+FCMAqCz9dJd73/JEQfooENETQvMMe
B4tiy0gqrsA5jEh2Ap02G2qR0zaUeXUlmp0kXjvjvuUV31xePV+13qmq2t+pkz/M1JMsutRH69CQ
8pWIY3JNsYfBbGi5RI2Hjl3SK5xLfl6KRExJ4SBdgcltyqhulWoIiscQLrk6dETpVWGCojtNdZwz
OYvNgiAIXeopvWd0x3+UXRxxS3WiiFHQo8+N5QVgJPh2GTWig0V/e0min7pZ1/5G04vCZc9mxRhm
f8P3fKDN0uqzDt6jv7cczS4WGt104EOiZgI+6gXt8A9uPi+yY8uxvYPhPFkht0ViMD0camEDP8Qx
6bbCHXXzd6fcM7CaRVhsvs97YmYRMgo+JgO9HvqlU5Miy7Cv6wBr7C+y4oMr5B6VwStkbAi3qsNG
vQn07MYvCxSNAQhHIeEL5QlSK8kIJfVwx3P2i4ueV0s07Vpf/3cAn153k70VFj6arKQgCmLx9aUn
zXMGoQbO11zlk2wHpIDsYNFEW2N3ta3HDu6OAQS5QMzuQJ6f7gJczjyzxhG7cVzQdkC1ezzcZ5aI
An8gur9U4EQhGgjg/qgTxksKZquh4Le7qRj/RaD7VvRcujfZfXsIOvMOR9PR0j373GXdtR54egba
mzn+35kNc8L9CgcAuDR6R4Cwqi8o0Badhl3x8KfR/Fxq8q3kjM9Owe56/Z/c35qPTnH4gxi7+JfQ
BHJK9SKGoHyYGhwmtHYX5fI6WCckx/dyXckOP8WlYJO7MDK3nH9kWsfU1WU0bg4GVZQDGvuF5lxM
BF23XIU8HnuhQgcomf/YUV45SjYHOyhMvNvH0FGSFF7VwoCwkjzhy9ymZEW9vPrVCNXZXbqigdh/
ShLWgLmZoklf4SO5RtNffPqMvKzvbVpCPBOxc9malrzWparbfAEDNMlLISRKe6EO9FmgOiE2bPHE
71RX2ElJ5wGZcNYPjJi2QMD/sDFo8rFDFXS1TTpIyinXyEL0f+0mUCP7MybJVsxvkPfCidfc4FJl
nLlOmp3vUW2hS/Y2IovQdSLIT3PaziZbjQ42DvAeriXGvQ+HvOhfY62s+il8bS6Jrz66KeHGNMTE
VRSFhuU3uo1/FCzim3uOe+vbz+keBpHDpb+sozDlEYgy2N47cZXLKct9Mr5cMvCToA5tYVAa/XLl
+Z56L9oOB3SQpYkoUgZ7OdyNtUgKKhq26mGhu0iwQBANDq7mSkKuwlEt96aHqohXT6jS3XXG2wQl
bl83CnFaKP1QaJ3HzljX/ALruFOkBPwnRpDeb+yGUzBcsStuAA7J4dRI6Lr3KB3N6ZInPnm+kHyx
ueWMvKsnF5SgrM2xvAx9jF9wxdAda+Bzgm05mz78gwMZOzDDCyCsnTpo8pMZDPC/afEP1gheDSFR
A7HonmFjCENLDmn07D4G5xEnr7QqtDDTyizfDNGVhetXc6bjN+9h5iprZRlCyHjuI/4H4lxPerHb
ARd5jT2oksw3KxmcB37jl19rG6ULkuGMyMfGLtlYa4ovRWT2RdN1mx5L3dO8/WlwNmC5iBrk98xo
O1cAlH3TKWVON36Xl4ibu59HLWUhgcIMZyVkEo+WfHVqoagdrszEdsgBmEHEFzjeEIZYe3i2bNce
2jHY4EldULn99wObblxmMwr4aZrFmZmTO3k9USAifJbGjLUDUesPbYr9yoD0W1Z9Z9CAyzpw4nOQ
IrDEwps+PAKEfCbHtfQ0Q99CNZWC1mDUF9eMNrQvheOzCAue2apU13tOME3kT1NWGlcWc5QqzR8r
PN0s8IMuwvIWfo6oVUO11Z9sZC5FqAJLJJRbsiUwP0UG7LBWr70dOplCm4AWl1jV2V4YYBin79rD
8rX+yNJqWAcy/qXOPNk0cnf385l2EVBp6hj7LE9RA/RYugyZwOE6zVlSqdsvZbOZRjKMUblAhPEh
qSODrBmcudtouh5Mo3gBiNCHzdUBRWCBrUHZoUxUTSnGdMCyyFVa5QZiVOwBRYchmaDLTY8T3pmd
I2x8ILepC3QxfHNwmnIuTf1dQvMtnLKloMVAyOAspDJvVy/c1E4SLgqAGUak2OwI+Q/XdOg15RxZ
3489cLsXw39Bh4EvXv5QefOGB5MpHSkpORoqGYFVkjLaTG7/Y0cLd6aq7IDcLCBIDeCnvM4qNfbl
lTi5YaBQPDiMWm2/vlE0w3roNwytSJsTgczPV5QL3kpddhY9k7f/aqvEigqrmCaJGL5SCjkGnqEr
TrE0JLxfl1DyOOn4wL+kwh5v6YKuAI66ZQ0jhgwMECn5iMt5e618kY+rgZnHAPAYSXwkbUywqxuh
bkbxMipcMvNuO8U9PguWPNS1+yqReLvIRCjEz4Wu1b1naUvbQWkQztD0nAf5OnEluub9715QvsKz
juVnAkg4NXXKaFDSaSwAoyNC3QCKque0C1coAj2dzezHoG6s01IH9ssRDQzOjHS5JLfgHwj87HMU
3FP45vNfeaZqRkI+6bBPK+tVN861PsrhQ+g/ncCuUAHCFSrWmXBiSGjzOyGYC+8eqhAibMr8T8+6
JTiEF7hIDqKiPIfGDJ6SNBjqsDkO6MJMnwN2aOmMqR60wEKd/MM0mQzokjfatNCdtWmdGSJ+0fjH
1xZgICAY73ujbt01EpnPprMp7ni8ryta2bnXFst+ZVzPu3RbQC3VEksPu1099AmxIaN1NKYYvMtV
1mevsKkwDR4uNYaw8ffKVunK/AMV9HJpd4FiOA1FqcOyTxzhoy1aUSRG2JTCRDhSIPApCcj//PIX
tsohuH53yicW1rKAVdw6qJmMrRKjm+REPu8dOrFVfLXrkmqTETMKQdCpe09DcIFDAgCTmy0KvNc3
WKOWoNFVxCrYwhE+d7YLSFauIfntjPwMSP8uMFxc3bgKqwvnhWSJV/SAuMtO13g3IBvfFUBct0MA
yGSOFhyJ0Ro/7tGjE+LQ19SB8I/vKvajTHcmDn6oQ+qkXpT9msoTzTLQlwy747aMlhwgxXgJ+My+
tQ8VX2xAVMYwIzEd6Xpqdw0WevtoLBeCTjWen/pPuL8wzFKLj+zbr/tN/JnwkDD1AuLdGIRyqPgL
HsvHsl6ZcirFCKwPZrVoEwf1WKmIXcaVkSuR9KhSXvTiYPbgHe+W/SNcrI6EV2X2m0D2m8j4plgM
J9E5yoP9N2zoqDFZSqEsufIRuFTJLZKmDvI+Bw9YBCzHYvgnqXuMHDvsezhKfqoJEUlqieDVUUzr
KQVzSMEfg95fUJ87xo66qaCXtznqrUyr24xM/koYIkJl1k139ifCMevqRgtquhu+Spphkpxkwmjn
JrWXTTEpnPL3wbaPjjESYUR9GlvtvBgBqbJPblYg8pfvY1S68xDfvk6CuBB3Ks+Yvdi3a7oH3Ylv
tWq8es7bl91Bpba+1yU9p9y3VPyJP4PuHHQQTZ3XIWnP5iMQpP8RkYBmYgj+C5lxOpDcozXinx+R
FiuJC/J7pCb6xBsj6o2+q8/3XcNt6UdjhOEejW+g3vmigXRseTpA9cx/3RqdG/Xg1hioOfjzZmS8
7KHOWj9Fb6hsVvC1RPP/k/wD/wWD6bszcDpJj4vg6iWM4L1oi9azSq9fgzziJuCbpybWdioav51d
x+cEiGrLbbjJm5h1eoQsUwRFLd8mYbYyo7Dq8DsPgmOpO3JpgXdtP7E4MA7gWU5mfWj6TljZ82Yv
E1iRvDszhs5UvBVled+VnZVGRuCseF34Ke0Gmn871b2C9HQNlav1WZkqKpxd/TL7LsePYbmJjrZ6
7ZhhmCTyBLsvgZiQEk9rO4E4JulcGKB+wvBWTrX85WZgQFahJsLAZfcKLYzrhYHe3CXJ+o8Hd+pp
eOOwJedzxuilFZ5g5X4HYHzzW1446UeoG2bYyGRuFhmE+XniZDWKMuSNP4IioMSD8lvYYXqcXoVo
kgUsGLtSsYHXj5hSKvioK+/hUukLNupUwsbx1wAYRnq/Yk0sP8etHKD9GuaEn+VpGsUxzDItDiaC
kOsdOs2cMbMf5xEpNfAh/EV4J1mid6JJ/l53DNZM4UPCH5bA1IisC5vCSEmUIigMklWqjHADpTbt
Qj78QFFqsH2A86xhxeZSXFhH4Q+ihOZQS1Lhi2Q6zrtwEL7MwMAPu7wPLUA2Eo6ll6GMiysSnDYg
hIOy2U5RpO9kJwNFEt9Jtj1tYr0tGmMMxa5iUmBk5gUS1ChGHXkseB7Df+Bq6mEEZSRGaV+0UgQy
kFvJxAYKSoaRMaDIQKrhnqBwAQaTwvgPlr+TGuMJ9F6Ifp0hkkupAfT4L67V/8+HCmITQDJadq6f
WfkCVytDuRakdTHvKFIkzTbnlCNqm+Di7PP+FROfGyq5QYfvo700QvBIynR0G+TtKPYRTN57IE67
ISDN/GGQOsCXalPAVABjHgK+0vaaoOCDeQAmG2eHQ23d5wXGxyRYvvNbz0b+1xD0Wy4UMbMswKLL
UQBtaV4I/5Tm6kUiFdfXtnxerxWNw54RQ/vqq5OJ7tVkIzlPIYjpwoR8LzN/+BltLk+lI2iexbJM
uvWludkWcLYiIkUmp/gTIdi3+tFPVOP3QxkNAlH3x9KwU4+tmUBqQu5dhTbi7xfoa/MsBfbPe40I
rns/jqlqY7Qd34tCVZvv2QbYzZsbFtkKRQTSbtvmdNNYC6AeUtiuEsg8pDPbFfivjPIcg550hdOQ
flFdeDBt40J/t7RpPalt28xouEE7RrvxGYOQz1lb1HlxOgshOVzMBREzkIJZBZrLRupKHwGeNBFQ
yngfz+2EP9rgX9JDUAvfGVGdThYSiRuJqRH59RbGM1K9HRGc7/LBnG82NWyvSM4EUguYCp4gqFp2
+qUUH5k0VGSY554rFa8Ls3BfRcQ/htCgg9WItxGGaBDKdB3wGN6R9XcarhJNRwSOvV8DqZ5TGsco
GydiA/2Rb0PzOetx/E88uBHOKlI3SeNHPvcRCF9hC3zYNM1fUQQPGafIAVl0eQp7j4YrKxzxIl3V
LXIsyQJ6zpHgIKmlq7fl2jKCIV65SYpR7iHSHmPj/uCQk4UBAKJ0AFYhneXN+bggQWB3hG2rLQei
jSYfX+PAiSe1CfdWGMiQ0/JH9Ogtpb0cg11AsNGKHdhRI273fsFueWoMTpgy+Mgju0ywoHyd2gOu
Mh9lPNjc2gr62oFecvBDPrfe8nZwp7QpkyZwhyyeS0zBKTEhoF2/J7n2h889aqqEryBQCfIcMkEh
CRQsy6JyL0LKRuv4qYOWTS2jxTVIkiX3UezVS5Ok91EJWljctOqVCFuJzT1lNW+j7DAASlEkJkLz
254LJbQjQ3TfH98xvtJa0YNh+uF1nngzvWIRm0xsQ5cjfHn95UFiHPUpoH0Qiomqtds1wiO5vRTh
nFGTL5ESB6zP5MDulgXCRrp3i2Zk4TWOApYw3ydeWg7AEDGyiY6a5y8s8ae/rr3+QcGFBsNO8ap1
5XZOLNWQB5DY7o36AJ+8Q7StFpqi2jQaMHZ8ERlrtP/OTdM/25eBCSdlXgjw7YHzrpdQUwAjXpAM
5zcEON8uIBRHXdEslnFdk1ODnOC/R09hlHYRahr1OJUpQ30ug2hb1yTAX+EBfRjMGlIg+zbO8mxh
bV8YKvf47paWyqmiyrKNcriepTeFTGjpodiSFfKyAHeIfMGQXwVsWH0gn3dOYXaht5XIxNcu+wdK
JD8MWwBp/nQSgBwYcbChFVtzHP38VpsB5Ymkidn+XMv7HXQ7BMeougmV22La+luV2Y85i+n6/2cc
sPZ4eoaOamGYKnX1QovBFy4LRjHHHFid5ptZzWh7wDkP1Zlpm2lCl62UqHjxlT/RDybS9Q5gDq4+
jkpz4Neell0vfoPpv22qo0QGQWGW4hjikMFGQSfxlzxZpW1rGF2KVGIxUbXSmkiP4ydSkY9u01xI
jaVqt8OsAxkFxCIFi4DKZ0Ua27srxh1GPXIMU2iU088r4qlluBAO4tp0bkMqY77pI3wttqXDsgWg
7lk7/4hRsdadYe0EsQJqG5R6KBiCVxHQPvPO4c/crl3APEWQAe5PQ0aIBhk4lBJ6EmJBmpQup46v
/GljwBvqsqs3zEHTZR96M/2b3PSglCw9pbq65hfqTupLHC5E7efT32xIy0ie5KoQWklVpb6XRfIJ
S6yZeblo8lT/ZrP76nV2ZP3ZPixpBlDMFZ2GKOq8OpG1tM9sGEW3cFJ9S6ziMS/pLAXlgHv+Uau3
4mbO8jJcg8WLNMArDlezAnxqIegT+nrebfTey7yCT+B842l41BJVPAzAU5/Gn6YSvogEiaUnxU3g
9AThYXurlLKVCnLtTNvz9W0ULeIsyzpAsM0ML18EMDdJmphS93VMsPQpKbT+T5vOLq9Xk/3vBHud
K1TPvKKyauPPCMcc7COU3X+Zamqddbhq6/VUb+FOFzr2HIJzeb66TQbCs4yQO68FHf/LKoiKsh5Y
0N9KN3OFlf9g/Q7y38+d3wEgvPeOfkmqdQdO+GVG9dOf9jfgAhxkOg677kX0sa2sUDyb5jdTyQeo
06fJEBe/IIPNuh5xaQnR/71py5k6mQbEIfNA7nP2rpRvo3BrhM8lNqx0UCSsnjZw8WHqDq5SxpI6
ao+6Buod3xjjD3F8vGCYOMXz+fxWV8WduDkl7gozGrZYEnZ5D0TkFTuriAwOJVRgqNJrVQEgI3Lq
0IxiVeEU+XQKl8PKIQB5739C4aVQoP+GAfU7iL+3s6TJeaOB2hjh7BT//tXEQpX1XDzKQt/8pSTA
aFSgfaKPdKXaZb5SuF6dhWZBwSrhfnQPgj0mn31NGte3QIUa1vrKHyfCdRRcEABewyG2eq1uYIrz
07++n7o0SL/JLa1D4HSAcmu1txAZTqxfeXckx1yDXa+pnE9g3xX8XgfEhzvd6JHBSG5gcjB7nEy9
jLcFzOPomA6TsaDEDlg1I/OvDeoDtk6LO/tKCOvNCbT0llr/UxaaKiNYkX4xiLA4acxSUQuZ6cGp
W0QsJsnNZXcdkPtUpRjMBEn1LNlnMjSXjDghXBU/VdyU+ONqwZA2LtlC1ehK0lPZC7YrPb8gAXVh
ga+7mLwsVS38rTrxi65kAVKtYK65rh78o3l7/kpU61bZ55TtUWTYAWNSjhz07hdRu7f1FM0RvDj5
3WexQMrqxE1gpUpjpYm8pxDx+lO6dcSsHCkqHLJn1KUHnUOki440nfA6AE/So3/M8AALc6s5xDEN
srEPSFr0isdTRgil0ArbYtly6xg2qikEkKdAtAiFBjWjtHOJ+Ro7okODhQBofYs2FJqpSFGv0JVj
L4VcqjSAK/CnHf/imMCS7ehRX2vwdz9fjhBeFbFTX15yLZoj484aWO54HFurvvMGpTFYPC+FOZPf
/JAzRC3yRTbftZydCcFPs4J1FHWxT88fGMxQ3enRZiSxYH2iDsXsAE4Qo9zDwAk9UGdIgArrxZ/a
fo8gYJE0cAEYOwEQwIIR/2eWSvwam2/BY9NBCdcw+I8jaQrD97NHhNpUcBeUe991m7xtqgc7Ji2p
61A1ENCZTkB6S54f4salZyFqaSo02J0l5g+1wkWsYnr4MMET+B6ZHCbxL9YVByVA+n6UsTZh1GdI
bzVVrMRloRSmUFrzEQaD06cM1dKwgjiUANTN8cAp9RtdI1aCvgTKhBgxBsdbtv1kyOPSnrWuJ8ql
mj2SFcZ/yvDb5ViyNUuSEekfIH1nYDMta/ydm5Ow3KDGpGa+5ilD0kYr0znsFNUYxusjRjjTXNVF
c9S/DxAFYWQ7amESPkknPULtMffeClq8PbBJ4DNe0SwaZV7PyFS/bDJNpwGAnROiLt7HZrCQvQ2y
xQ1/pGu7anCOAew8g5t8BsqJLYPGsoZsXoktce+2ohzmdfKkHoV91+w9hijdlYFPKip5E00/Rc32
veTjA7ey3Db3Vzb0ncRnH9EplDVdf/G7h6aiuR/wa+0VL+8MlbA+yCWO9FXzrSAIDi1qN/y8B+Ra
+BVO5CWIF0c88QR5keBVSmV1ItX/AwsAYNgvN1sjdRvRF2M2PKvyC7jw2R835wT6EWRzD+KQLrbm
3Y29EGHBYnfU0bDVVf8rXAn5p/3XPL0TGFQfeCe0UFd+RVS86SrZOm6nbLuTBk8AA2Jxjbcy7vRv
pjU1Dn1fdR7N1tHAhokJ8xMowL8GWPvTiGw+yhiZzNRVKUmx0rq1F6fUZ7akv5uP7lFBrT2RbwOX
FxQy9gJy3saYYkZR8+RGy+uzTFxrK2Qwe/xbYBO+RSrSVKZp+uqFq7RKR2ZW0IqSkPCY8T1mgU8y
tB2Js2PE/NzsCehWRaGnatATpks2xU86qcSXDCFn0qcpDN6PWsSePA4EsSdBJu0qhQqIQFYujMez
8OKvwEzW0m9ZBHM1rLOW5S047nMuvPNvJxFPKlfhu6HyantGaqu7SCCxzdxqxXEmEBse/D9WTzmz
HMjGQO/hxMq1uCpSB4xzdWl3yMKJupIm1wcd9L+mKhVpIXa+fdBJhdqouF/1392+No0Ap+gy/ikm
r0cvn1y9UlqKuozOyviCNuRxaLzT9kZ7zcWdCTeFbdrgWgkTBMr+iOkIue/6pEUmpQDQYW0CRnAw
L+MASAYnuROof4dqpw4y7iJROcEgmFGVThOfp5efurLFKyBhbunozwZzOeJnZGLN6iR4BVd0GJSe
OfQXLxzi+OFjMuaSm2+qHRfANVgNeak7CFqXLsK4n5zIUX4FmQ8/NNvE4eAKcfw7p3awnLYnQPqx
WnYg185fva23u4NQG40Ok9pdaW+8svTqH+iRfA86TXz55P2UcIru58RCPJ0n9ZDSlJciQRzbimqx
p/i+qvLkgpN6tQScsP0yJSrNy/bM65KSBZy1Ur8i3txBB9ExibVMMG+nNUjYlqG1begIkuRk2cKe
IonTkIRh0abGafKvmRqSqUUrv90BP0JYsSdeLJJmFq4MRE0elY4gbcpFJ1qXVuf4mVbXUZBK2jF8
IsyC5cnw4yD92O2oLDUgTkv7stNJz+QIFgdziaGM2M6bA+Qhy0ZTdZiB0hqjnjpcsUY9+XjSjkMQ
8hsjvPdC5gvPPNFWWJ+zQRPH01C5H/dXDF0dzKBdJtsj/ORB2zK45RkakH+xWfuZwYiX9FJ5AB+T
Ai8RoZHJ0JR/nbri9KikrrD/s9m8Wpp0hXwlWbXZQFALIFfJcbHsiy7yd+EH+cwiAaRWiDxCeJyu
/RzMzgij5YLvB0zqSEWtBMbT16stVLXIfYWvVRd1Ly2Xp/9YbgT8wIG4/Zh8uV6+6bDszyGFOuCe
Sc4173cDWfB0Dy6XLFC1LJlrBVQlR0neZr0hqtEYYAdSYnPldGQB2GUnrBz+5xGWfhBAz91zZ+4V
30klD9flk4JccRbXHYTMPq4pIzrMFHr6BQ3ZUjNpepqWiiX1AHmrWwDQccH/ZE1lKdVyniAWlz7g
//L/3EifWgCghD0u7RcctAKhSowNA8oVZkWtSyr+coljKoHYh1D6PZD4X9r9CETvolWaEPx4HFuS
2rPqhoCEBijcRcAauiNW+A28JhRXKD7yehQlU6Wz9BFo+uVP73Lcu/wIc/AAbFJWGmft94L8PLqr
7vGZJMAIzWdKMAJvCxQRdoaFhXnvIt7z4JYPqL5q4kCk5E1QnLFujR0sM6aJ0q+GGCgiZpkSyIL5
nXUCXtCm/SwVWYls/dUkJ4/hQtZDssszc2dohtTO7R8fnPzjULO/y7C4JKNXeRitJVnHBFS3Fs4t
OY1oPstkOmD877K9AdN+BSHLVQxh3uy5+SZNT16BZFWOSmnvEA/YRqASpR4nB/uziaQb+Ilk9FPN
uQOWYWQzYKCwjFPOKSRkYl2kt85s2iiiyd5soBRKpt++OQTZl/v9UhJ0LCQCuamOZ1hnYtu2vjyZ
1khQWsmubGXrvaUBl7jzuN86e1MrPTm9yC6XUtDXUgBGS/Ij+mg5Bx0jT7iRAaARQMXAHA65mbMm
du6h+EMJ2oArl2fcd4SgJ9rK/g6+oPiLOlFjWcIOpCWLdWQoXG2zOoOH8M95jmDqGkwG82uU49Ne
PvXIPcnfm4WEjeGW9LTO854dS0YVcymwY8IYmm7BQwGWr5qUaxA9LdObD3zvOrFMbSuj7jB5sobb
j2X23oKz2221GErWi501m3yFle3E3/tRFT6Hz+59S+wM3RK3jeSiOU2LPHYIQ2R4JfQBbAnw/oqI
GvBF5eTKQbUpBlsX0EjFrdz6GvYpe0Jyk6BUojldWAFM172Uwx0XzkpGGuCKTQA4Wrm8jEpOo9I6
qLe79yL2vlbBF8Ov35fIDhxmpp7ufEcXv0DpEDoY5swMsnHTPaFQc/x6je03GlqcRsdHWFuRR1Jg
7ZogPCSSmhKWtaRZm09YGONsHuLPA+wFsKRI51Kxi8WOlNO3R2nlPK6i1NfeT26N/AHeGI/MzYIE
fNmOonvtkqecwPkv1ZI4Svdl6BZtkkatZmxHKQ9eGLdJLGydjqupDQYn15Vo6PHUrsJ3Rl9vL/9k
TEzTp6f7J28y7xF6pJVGmrsMhrSt3gVPF7phOpuPoZUOm6c8Ijxa09fd2lk8bfjuFf6mUFzdF38v
PcVli5p088U2bQkhkNDM0opzZitB5ecC8geiTaE5EijPyxO3f4iddyQsmGSGgLkSvswHCEzFVrvY
Ja359D9Xef5g5rXrqgJ1dAoOh29l++RNGwtuU18NMZn0rI6GESSWixtIxEpdJd9w4o3CBsIB2f8H
gPXtQpTYGYaDZnX4NIIro42HlqcuVqt02ajuq6wIMDyRyHgBiC3+gc4NOV86u53Vw04PIQdeSM+j
8NrtjOGTiHKooLJIqIL3FsKqTQ9+N+ZuQy93f9KiyOAjPS27Y6tNYnhynlSfUWDrREA0hd0fngMV
FTmoeZ5Iaeo/Y1qdaYuk42tPziuJxozfpPUcATXvehvc9AhsYSavdyxhz9fEYt1U/wX/3Lq81RhL
l6TnmJCgByhd0qtMjfWiK4JJE4hj79ZAs2x/J1HB/JuSvGgGJ1j5O7YMOJaW5fl4jfaE3TsvEJfz
HWW9vHAqw3QCotYor9zSd7oFZjjUY2K6DBI55Wmr/2XHEDXSk1qThl8iUocqF0IjKNr7An1JS3fe
JRO+nbQz/U0no4GUCPpqWEkp1VN8bPnZHYVIJ4z6PtHuuF7a62YhXI7AfoV8IfF3mWUoJxomPhld
wLgNxij4fwuOYWCXNiXkxGN+f5cOVmWN3DdFaSUjk/YhetO3NLEXUWyvilXBTPfS4tj3ttLuKtV1
zwrLdQH9wfomHvuc7UT1wmwD7x7fxV8La1Go5JEL9XQZRpvDpBamNPBTKXs3+cU7E4HKFEKCy4kQ
7n1ZNZmiLKJNznL1e7xVC+ijwuFpQ41SSdqsHSYF3aMgRI/CfYbaLu+Ld4p+9DYYv16+3MYA8Epz
pzePExiNmXXnmkv7+XqqB1z1OrMOh5LF2v1NVIMVxASJW9jJf50WlklNQXjMfh0v5vbyvQkZU84q
WSOzOBhmsEi8yxbveHeZvK+jos3AYqogqXcRPc0ptxUbuBWDuFsqs07Y7fAmV/fKjlDLYR7OtjAH
jjP0iuHCWsFN9p7fm4ckkU6LWs3XqxkhHNYuq9V0/ns5l8cdqgMK1HrWKmAIjkdnpxB1CgSt+Klw
C2G/rGhGp9md6nWtH4lip7foDFL1ZNEcSwEAILEgSE8MPpwVgU8npiGxpd1K/QMkRhnb5oJxoVCh
rt/lT61gkBRiv4Jx+ZfwemAvAq0RzgE/KYCXfmpQ+2vWR3OrApbFUuW75/7kXmwU1oIIFuAaYm9A
GRnCUAd2DFOOZrB8RUIaUK1WjIMafevvHQyKnZ9fuFhCn+CjOQV5R5t1x4zDC7ZtBU97JTMl0D/I
5dVw8Z2j1MuuXTbnMhDEi0P+Y5+03z2qAEJCSaZOzbVtuYsYM8wqILyslZnRryd2OBBpOo3y8b2X
jIvRd7aCOY//5UTxJsTKPb35lXZ9/UKP5cJ3Y9iq/k3F/tsBlliYgO60DBMamj/XshFOqLPdWWrj
srYDKtHN7PQWwEuvwQdQYTj8PZarZgScbDxRQiYDwRM3QBy/Ez0b4G223wUOEjxb8ecZFgYFJIKb
HTGPZisqttiLU16mvpzsNicyYRTKw2HndKStEL1Fmkt49Khy9RRISpB4byygmuarCOGssMyNcTAJ
JMgSGIC2+8LNd1QX22dYQC7MQtpsw6SrWj2sMbdy/uSdJuogKd1c9Dd/4aIuTJ8nRJVh3e4Z5a6o
udvAA/3Fr/zBe4l4NxPdsRfDXe2PfwE14HzVGY0zwm+OJ4JRo517l6F7NJQ9Vn3T+b5uep9P5H4L
XICyKdmzLl3DCWgPfnull3L2snYr/2dz0IesCXFq8Pb7PsJHc9eiuDge0bwRTpLDHMayijGVKg6v
UBjhfLSmizFcDCag9FW7nsTMash47sOCOaPsBpyZnMVJF4moU2jEGpoUZ7gqDjt2AtNSsmkVq1u+
fIoARBNZliABrCOqNQHhcgFh1YuJ6ZEsP9+9ykV8mhyWMl3kUZegDD40nGTLrtwfBNJ/RgWshFq5
IHRvwWP8PuE7oNU6MocONQ3qTNtDTBz0//pD3M8IrxDZvkrQ8ZTxYy4pbCmA4Hb+EIx2CzxOlYH6
l7ndtGyrO4aShlAcy8Mk4DJahwh7LanLVninU5Pr/tuT+zqmJahpXA5xr+zTJTL7dUzZmvulcRtX
gAxZowtvXd+MaJUL1enpJB1wzdaduLZEBqTjmYFpo57sYUOahQfl8GJdCfRIrsOGeVwMM5kp9lH4
F9mt3bo8IJeWEah4uyp/J54XuvgoHf+dt0XfeoqTKjUqIzZO1FgzWNW8QX6+bOTBbG+HG7UpaZg3
xoprdeacVh1DN8GVtQaDK5NaNzz+uCVcX5Br4HoZeeSJu3UCuARYsSfBPG2d1S1k1LtqjHHMbRpH
vz5oKTlItNtKrb/5+lNPg7KUum/PBldeHBeMhsc/iN9mqhNbAHKgep8E+gYevCau9IhCkIZpfjyj
3UogxoBW488SbBKTC+vLBRr0YT0U+yo2xxU+9hP3hygjdnPgvEw2V6lrDVSKVdu/vRKozZfQL3ql
5qa50zpTMV7Mvrj7JWG42IjodwAV09dfYzYS481yJd+W81qRht89h0ZTVgiMALA90Uz7O2+S6VCk
U4JCTi2gJ7LCA/rVgIw/4tvPDolNv8m59pmlYgMfhC+ulw8VGEINcsR6ms42I0UPJA73VInNmYhH
bXCJnP+6UlBs7oUJGBTGg+Umc3zd3T4cY6K2H+vQp04t6CPNtsQdMF58lPbJd5uxsEcm9D+0Xr+z
9JPqFEoJ9pPnmf+rxa7Bi8zkX/Zf+ookMKQ354G2d26l2ykbFoHk/GQUTvbxwoh63EW8Gebdf+Dn
UYiDMA8wgl7O29B8nEr6OKNsr644BZIn7cslqOvlDJ0tt9dK5R+KiHqPU61X5pZ/eQkJFBIxVoGd
P80syBXTb+mc/SnhsQdiRT0ZTt5KwVQHFHRvJEQsqGOMm/NOl0qqmaGonD3AF7NCdTO2Gtl4OUZH
Snk2JdD4bLOw7g5P376WbD7JBYz7AtBtk9u7fgNbFdHY+5hJMtaw/UcMOcb31zVo70v+2NZh6yKO
BP3+kxvaLfYUGclLGLEpDkcvMYV5Ub6DcXw4/rh0OR5QqlJBqeUmZBPY5tynnkqLAoX2vt3B1fVC
WKijkM1VS61btA9pONoOYcSRea786urUL2LSOM2/C6vuRoxtpx5LM6cIK29LOjf7KPeQ2Zb33Nn0
V0JEHb9iSFERdAvHzfgvrn8suLH4LWFzRV16x3M6OPqtohzDkQ5u17cPkh8fJ3Z+OUkMDzCIZL+k
epMozxjNzKdisMUi4NCv9DzlfzslTiJNgXkvbzJYWbKt61Ihh8X5AyU3qZqKJuay6wQsNVu7q3gm
NEtfAAkWzpmesokzEaC99G8uP1WZvnF7/GVjV9r81eIx+dAqUcr93Cy01TQ4Bqvn1byXOc4FFk/F
YkQuHvmwbYHehYPnXtoU6soFekzI4csgwzilcAXMAOTQr1dyRN0Ujz3SYptfgt+yVklLBQNtwiF5
LTL1D0UOQKDv1vCiNAO1b0sMkK6SreZqDuGEWBInV+oH/mMUWj6VKes4lseiDIBurrHPM5ebnUm1
MppgUQqL38AQTpB5pl0eKl7FqrVLcAjZtrnOkLelDCGRkQO/CFIQ1Jf4xrBADVS5aq70F4kbWo0W
35Xu4QxkSj2EKTLr+tRllgjaR8KCq/fipnG1Mo/RwmtOtpP+YbnNxTgGNm1QHw9CYaxvgyTXiNRO
OYL3wZywGIhG5LER0R21HQwrXTjYuPL3vRKDKuCjCmCrE7w4oJf6xSylDPrEtlqpva7uHLdgqPs3
n+9UOSX2/+LEI3UoqyJ1Hlb94KvBIaI2/88nr4XdHjomMjocYifrvOd2B5H1n7ohlygVZ9ytNeSx
+zQ08ndWphI2Bqx/WBkkCeki0DZv+ovYx7EnkdoM9z7NR5ylhawVlAPHctfhwKJMpFuP42J+Kc52
Wn0P6S8dcg/B7+OkG8bqJb9jbecJFGHXF9BzsGSjC91yefhTrYtn1YlZVkLRRBhf7xJf+U3Jc5/o
3p5mS0TyFJrp8L1Q/FTNMk++++0RuLHABguGycGlMOSQVOBspXJoS5c5UwCgbm4TD8t/RR9VHxBy
3mkuhj4IvjYaFIw3DlidSlM2YWo+dwqdzbOkfSi+MICHvTvXgAAIjUhep5xBCoMpuuAOqHy6JqFW
j4w2kmjBRoP/paGtXL4Xea89GEW49sFCUDniaWThxcmwLydN5eXvZRMPAp6WLme1I02eptMbiv6a
AccnKl5YgOgDKm58nXeS/oGj1aLNHSV7pDCyyVt4CTO8xitlmJlrYDhY/ThRCGfAaTPdpP7lW4pH
4ucu8DRl2fZ1qSGA2C6fdEOTbya3DXBbKd2EvIIuDewGcWGxdtLUHqGnBq4ijC+7yRB4JU/qN2gd
8ZYK0CtBHJVRqZM+buAYx58A1VNSziE9uu9E8Zo/2DCG7WJFT7IPqqfFzVn3Ap2v3PVQa9MyoGaO
1p2COuyylUiCnTuNrhitg3eXeZwGYkEvmbJU3tjOjkvcQzqQuk6AeLFfAPm0L5BO1Xbis/4goJ4i
O6uo7qWW+hyialh6bPA13mkwJniUgokga9ur19U6O3uZ2yUlaB3wRFs7fc/cNZnUh/fkiQHXDY3P
VyvMgTIzFwF5F9nD3L6YWauGnRXT+P2JytaNzgL6xOWSQ7WU05MFylxGuSSY1feeSIxdzmjHbmha
EHOS05pRQya9kEDPImbQI4XodTgvQzoV8VZvJdwJBXx2Uwn+GOnVCForRcpajLmzjhHk78qdp33f
OidIE3Nv1LnYcJIQxEU0YVIWcdWQJjK/g1kgziDD3Aq9AZv35GzptWSdAn6EJrWCUlvNEOoKimFQ
OBLUm5XpbziRCUNzTi8hNrTeSXvSp5s8m8BfKBBFc227sRHrBrHcnhWQb+ELhqt14VglUrFQXB+G
ZEF+SrnsWJAc1t2Mebsf+ddwyLKE84E10fGSJG7uVJZOebx6/3bbLHfxcv4BAAXUHyfNvSdfV3Zf
sDWOMSdxeis5t1wHiag0yCs8BSLQ+DNtLXGcbUFS4ctA9/1cx/zE48jmohbY3mJlL7SU8uPQajRt
BezEyUmq8gaoEHqdiBurQuzTNt8KtVnBx7wtcwwR9rMPnbhXCtXXAihNLBNakECshzubwuXQP8nF
K+H6c91s2xY25sP+BLXlB3xTbAlWegtOfngCY6KM0LwHVBk66eYu07iUS2z8Um4sWs0XMdVllPw1
Afr8oQik5CHhpYsuAYWjylP2kbKI3fjk4fClw/SAw1WRPkfBRrq2W1ZwmQAw4AtvLEw0QIK8/89z
UmG4NNSD+9p3pea1UFwFo27QwtVX89PjLanZndHxg7XFwokGtegdisuLRLJvIT70fdO4YbKz/8da
7UsazjT26WAndde6bzdLzvjSaT5wuapEGEI1ZMCAK6JDXIiCwFaRHKq4jP84wLGVxk9x/9XyzRFx
7qDypsD8ebz7tGjJaz+djLa23I+z8f5+ztlzNq7yp4FZgsgFw9tiUQibfxnzWKvvZTKwcmEqSd1c
cMUk9Xwa2Iw71GQRhJ3YKGQOIgMDD1OUh0C5nlyVe6G664jfDLTuuzPoyPTqTCBqdeA7QagyYbgK
WXmHWxSRtcCPhC/OKiJQlhc2gaaJPYluP5iDkEjnpNF9pUGDTc5rpdLo3MEi4qwoXcaeFUuN73E0
hnIbsOrwuM+vrG5NHx4bso2d8Pv/zvqTj9dChPUi8Ejwv21Va1+qvP9luqbublBJ+vEJ8hQJy3zu
K68FP2tq6G7J2PqiXgXVVxJ6X3RdiRFiiOgtKUhbHhj8X4eauviuXyn7LYcKMXsf6wVnmY19wjU7
Nq7m34TehLOXvO6oSgFx+5zH+5uYjglEHcA1YOtn3uChBLxOJmyP3bQ2siIURfGC7kIJc3I0uAfh
/QC562ym6XQy8IUe7WDYsj/1douvm3jddf4r2i7ZgkKENImmqBSw5qJSFWmwNCx3mpfsSofe8Gus
N1kgvgdfNu0dTzBCluG7SmhQ5BiRAny9UGXUsERbgeqW2nrHDy3iln1qWvsv0L6O2ViuV49N+Eom
BVDUutU3S3RAn23gzYA4pvGbEsqA8Rtjhws+5WzwlU6uXPzUKhmF44FPHo/Lmk0Fr9qGW3P614yn
oNG6aB7QWV/AmYaRF1NwlinsDVeQkWVHb0U3drmfvd7VKuRZBISPk+Aj7YP6qduSL1QjxzEgn82S
sZFBpdwUZ/x4/oKR0JtK7wrGcjDwQ+L5vjDwgSEf//bQTpY+Zz1zF5THUaryEkDTzPV+AEzBsVyI
D9AruZkYBwnSsZBXP49V7q119wbEhtHOCBcRwIaC62Qk9Xwc+a6mEBjViny/gs0uIyWd2nXSvX4H
9rgeEYMc/k8nXYgP84hyCQUOrIifZz+12zuPbxWMAdG9swgqgXF5AY0hqfAgHIJ5ez5fLAunRdcI
RhqCuN7ABz5kM3eKUOpukdsgRWg4kR38Ds2vfK9eFKwrXqe2zjkT852UXMEgfh6L/OVQ+6A5yd+H
BgN9HSDDtmS3mZnwIldFqtBpsCWAXXpGUqV2muasCA9lKb6niWuRL+wnio48YWcVzctAzlZc+6TW
zGLp7whD+ATKilzVhRX5FLDH0c0s01VNDTFDvfDH0AY8w7n173pH7UsWd2bhbK1r2bf3hxq3Nz9f
YZW/IxxZOupweGafiemA7wclenuO8kAYnC265kN5dq0jWTb2E+F3ID49qoYFLeXflK1Dl5RQwTHp
fp7QPknOEvW+YwCLtY55tYirmOnngyQ6vP9pwtI6aM9CfAorI6F7Pzb1Zw7XXfsySzBvY57sCvy2
wPqtdE3IeTvAsspXzoConUKMXBb2DXhAgiGAfLH8XnJtRNgeRdJoe0/d0gsomPp96zeFIuFhEvgL
LFuyXrnKroWqNSTbSjhO1iIL0sp/ni61xHvDKW34VDk1m1mGl7yWCCB1mDRfzN96mrz8a5Vn33Rp
QL7a69r3zM7LTwQHI9fZdejhQc7NCx88mD5Zpd8qXDEJoGIllU8wEDOdT0PuN4tg+FIbmwSW2Hu2
69/byORdsT6rpfJUkeWmCppGrDh575slRQ8k0QvHw/nIQCtR5lIvBBeIJ2tp+btPZqrH+TtsMRXj
KCzd6A8t2vtQE9cKDUHJQbRRQz+3jY9LTaxhIidV9/GghxiChjQwTcHLkCxALCHbjUx0ntLPg9r7
V5BbUXV5JGnlHlh/nuZ/JgIUza1Cs5vae+5AbLuepsSs9aWzHpu3H0LP1IIPmgcfhM+QdY59dejA
98ODL7zA02uxdCpGrapW1hsItZ4mQigDjhNoVd0hG/q7Qk1qzwXbVKIlEBld1mxXiTWvo+S2kTM+
mrvuGX1MA3I5Fab5+BRIhLgMZC67SCEu2IqLXJEWtl5nzgtFFHNfkSivH1ffvlDv2IjglJRhdzcg
Ao2Nd/GPmnOCNDxGygu43/j4Kg2AMKZTGCusdaoS0J3Ju/xBs9japJ5A6uMXBZ6CE24zpFdLtViQ
KAl32/H1DZGvLgBxGA8ZFQZqexTSYDHLLBKiYn2x7nuPzPyyki3y5xPB8Mdq+/tzBwet6x1k7u5p
G7sRpF8ZxYpaaigBZrJA0vzCd7r0A7fUi6y8dvWksIae6k295eOx3oER/yhNEQNDlYYEpYtd/Gt4
a6St8sQf/+5KZZENU/dfLGTMZGUGina/+XPEMXbPdGDzWcGGQHbZS4O+/n2JzrbcgFY6T0Lvgjwy
8vbg1MkZIjD+yuvmXMsVnPVMPy53PYcGGwYC87ltOhHlXkw7AYHJ5ZLKjWpOwO7XHslQQ3i4ofkd
SaC5XmKp3jM+ncmLims1ZN3LrTAnAMxm5g3Min1Oo/RzJfrsf9aQZvJau55IrJc5UbPcpvXm18KF
b+23/2k0msZzG4l6o8xmwKeP3+hXza/jqwL8ShTTckE2h89x7chX+0MmvHV29SjDONUAmcNLdzND
nnqOmuBDXdPLStJ92idra3npTcZR0C/NLJ1kSQu7gvLt7o6bMBsUO5iYzKWUh1+U8SotL9jdvLZ5
dBcy2pt0NW5gWcNR8Bb5CBia5VuPtuhOboH7t2fU4KkrUEN4jJEtbIckpe+F5qDrYTvJ/btcOhzm
ry3513fGGVDR99Xav1y43BG6B3hI4asWnKbKS3VzuhYFi0r4AHo2eDpzri1Qa4UpjkXopD8aAD1d
ove4updR7a2yL09Kk/0cVpGhgqpBACE8ZW6Vvg4TTWpl2bLiGVw7ECYChSSkSD35/47UgSoio/Vc
7XqQrv8SEKPzg5jS+A3rA75/O7wMp4IQCXG1yVUB9v1hZ2igH6tQ+wLj2RdzrTrKl1n/sgcbe8tw
Mx68VkUVJx+gbvSZ55uKw623znL/mKo2d/+1JpQnOLGZW+gndGAKljwPsG3jhFcRuEfzTcXyIv1B
y9UiVpVto7w1RpYDqm/z6kwgdlVPIYNP6wz0w3wjai0KWYYKUmYFrUfP9oVfSG4LxzOnAHdCqUcn
FPAb6txZoqfOy3akzNoZn9nKRBzku+QpKBt7+gppoGlMBCMiiecQy8mhFDaLKh5TF2RNHIz2m/DN
HMuK2jiVNUiJ7Csuk56scQTBf+lxEZLjLVrZ+3RcukT6e6ITwoQXqPXBTpCZ/Md23HHHzvk190O1
QpqtqGhzXhozQh1WUKFDvoYiScbsspZXr16LtoF7UEaCudccl3rXtuB6TSbBEzVj6DxZUk0sVbdh
ILe0jh2w8Vf0LRgqkeLahW0PfLovsYodNqr5HEiFGGtzj7kwowbtI3seU8/mxvXWHgn3WXemPoEw
kgDk4mXuOSz7s39gcyGXkDYZS6iyrshYulbiDZVRIiQkXQqMLjgqK4FFMIQN8BqEarbJmnvlT18W
4ylhqKFHBV/iHcdW1c4cileh/Nq76neL8O3C7V2Awh5LJDbQUa3Ni2OwVKqIV5iUF5ErQUDj+1tg
qHSvCb788bstLP8UAOapLkoMRXWIXh84Z81gxPUolAAvXY7S+tCfjF6/lkSYjhw+4e+xda+o+gAd
1yyx8XutszaYX/vJBLxD3B/8+ejwyq+hUX9GLT6dN/LDittzX4LDkkSPHtfsCDwUkavRU4/vQSij
iYYtGcrFrr6g4QFMXtDMRLYlt4Mepzho12l+3gxAs8A351FCbDmwR3SLebkn75Ic/o11csrIVlAI
qEgQw0Q02FCYJxOgOfoJpdncZgh4bXohKo9GJo+NLhSY7HPW6XWTzjNgG9BWY2BHu7vTsH64o3D1
cXtDoj2DEDyP4rrazaA01+D11/qTp6itjue7HgLj6YR8sfb9vnU6xDYnylm450FU1BV7jeqHrEeR
YLnDANcsIGuVgawbsy3EX8xQtPUwTGIY1V+SiUK6oePMrcczu60lC9Ah2ue3TfcMyA3KeZemJdkk
1oWr3uigXdHy18ha19VSimoA9EBBZ/JH8Z/JEN4F7KnJz7J2drTlH/bZCeajPALxGk7nuS6vrdY3
JxTZbXd3997kv8eiV0tNCGpeAZgxx3M0aBWJFNj+doPLp6Zm+naNM5jMHjuyRkQqzhYNywoiPVkO
y9bJ27pfioLdtvsGaHIHsxCtKU3W4WOr8iZw6Lp++jp8i08nrFqGoK8UYNVJwMa1WvRXNJY5++bC
4wHEriVC9hVRqOI5R+S4TpLepgO6JaQR/bzls1TMEGN7fZVvcY+3bDTwiZWgenj7GYPcSdaHVIS2
8vofrOvnTTIi3D+O88pqctyUQ2DTiK5wuJhL8BcNlC9tapsKsOztbrBOe3adz5u1ts6JnOtZTFgH
W1FoEDd9R1aXJ8NuPjRkKlQou9HAvWj/+VIrHXwjet+EoQ3rR8LGNtjs5T4rNxLC87EtXovdgFCE
FSZbf9K7/Q23+D2JlOQIp5VUZ0D6UFLFS6kAZ2GOWFdaIfT3FvUXHjsNRdGD7B0Y9HoaF1V/HmyK
W/rPYh/Lgo/XvJLI51IuRPB4UvZBccDGEJmicWJ9kZIqaSMF2I6vrHZ7n3qzn8bfARcSf/mi/+j4
6Rf4KxvhM895paOrP9ioG5uhtgF3B9qcWFSwOaHDWVIoqdOddWe6m/g18vDQryeXr/5IOdF7pLpD
9FAxo1o86WlQT9eJSRp7wgCUi9OECYGcoYRFF5B/j1FcdRUt3bOMzBS6krODw/aE64GS+txYmDv2
ih8wtj8RJ/JuZn3yx/P831RMGZRvEQhVSQkzUH/l6DNkVh2Up7QzUyUHeA1dpA9uHVBH8BrQKGwr
fUT0kd+1A1gvLoIdh/0CoeCI5zEUFcF1lfyDiq4F8t1dxRGLb80rC1GDKWC7wcW5Fdk9f0HTKMOz
fe8OosgYPZDfpA1kJo9q0nf8Yc48IECRIx+sZep0H1jYFQ+D8ImjcI8kWXV9wBKoJMHHP+bbP+mu
IGN84gS+g2dUbwosQ38WHuRsoFk0leX/JwKQ1zR+MezeEZJ8cPedYLhZRez/CJkHPGtuKZEElsGt
WOb+uHyzQhLGNuO2sPfJS5PObI2Lc/nx2asrnaJ+2c1M7cSR1iGtZH32sPuRKOveI+IXk3iM8X0E
jVi+yXkh6eQJ5pPoUNko4vneJCDRrrW4totmqJQUpYnEitW/ryHYRLHZft63of6HlJ4iWMon5Yil
dABna3BA/pmIkUhFMvi1bHsIDQYK6W72fk6slSE3Q35L7i7cCW2NJhsxJH1J8q45WVr2U5qx6u1x
L6ekM+s5uzwcpvX/gc4UDS2qpvzyfmhwk9O8qe5oGVlzGOxdD6X1EmfDI4M9IZSAGw3+ePgMHNBt
14i+1pkP3vB29qPD7OKmiZD5O18hJ8XyRD+4fyUPEXs7eDv1M+hO6dSk01DJTsWS+coqMPRwFYzM
ppxJB+gscYzBAFQucjiCHsHybcgPvodGeTPDICpnEaaXWZryN3Cxf3FbWSA2LRmPCaFa7+/m2/pW
WKhGMbfhQb1DY8YUx+NXEuhyGO8CaUFjs2RrJwXv2W0Gj9uIcCbfy2Cyn0a+r7J2uDlJVmSsRXth
nQLF6dLo+hPzvZdOhaaZbacKI103zKo6Etf6BBzFdIRGZhn3/pqCkDa62UqNGXW7Rx5xAlvi5fxc
5F1bBJ07G32Zms5oMhFiOL9n/WAzGDFBOVrDDYJl9uqz4FqV1gq+B06Ks2djRWE7yT6IzEcg4gtq
83xQPKUSq6cY78Wc2qe/512KGYHkuJs97ttd7yG/mIINNJnz87z0tulD4RL43v2YaGVMdOwS5nS6
WFjmVd90ig6hhUs2OnOUfjIl2fb6oPn5ztm69ZHvg6katPBCNNqtDOnn2s9F8I+eORe7fS/wO5Es
IR3YOKC6DF7t7IRk+9jlY1FOLMIsvbZG4wh2ZsDvNlX8DA2Rz7nTdHbA7jIvFeXa/ixps7MF4CpP
a+I/EIUgHiQVl3/4UfourQpC+7Y6W8397mGJamWCw/4+XZGzltszKxH4vDmtPNL0hGm23LSYHFPU
H1e4VS13mKlI+jUtSCRQ6Bm45kWh67Hi1jHj4avy/qKRpJZQbjmpP71+pm6xWYS4mkBHQo4V2yQv
OMUgUwXOIz3TJtqZRZAw0GkBksYOAEhhGsCMGgDVJP8UH96s7uImL0GY/Vu89yv7JF770XBEczQi
Fm/HOt2zuSm2cZnYJXaP0Ef2B6UhFIVll/RdgwW0IdSTkV2NLk83EJYPspTpZXFNbPkgGBUJNudO
LVty2e1+G5oqX9C6R+y6CjWgtIIjt5sAHFdomYdDTw3LyJG78+BAA23cLZctlx4MwZBOw9zwVDtp
DhdymNYK+oaTsSYKtYZPFIHYWU8GbLDZhMb7HGZXtY0DnUjdMci0MrPdVg1eg61HiC6vodOnyB0w
uFdkAHvCqvj90BTXUa5KVwNqNrnluSS/ElE92ec+wqEETjOdxMTlkf7HLkxMBEgHIfd07R6Nm9dz
+EUQkDL/wXKxt/Hi0QO7/W6eGTP4FoEXXUDohuHVScXSuRH3vGscx9zXsQQJisux5oHy7V90MH6k
vbFgz/yAeZsPjYRfgXi4L/GM+EsM8tV+a+dheBPvOSS/QY39bmB01ZOa4fAiHxzNArLnLku18hIW
Bb2Nzmv62P7qzDH3ONJT/4ZaA+y9PkK5MHVrVxmYUVvuWFSDp2VS+Tq+VxkMAZcFNbEiNgstipPo
/SQkT23QVJGAwc/vK5AFjsvWB1ITSENzcXVJUBbJqRaE4HqI1mCF5l08NMxeyJijv2bCpAJ8Ks4u
wgmQqn+9L/E14UivJ1DWAKvEzgP2GTYmE8uQ9hIW3oZ6wQ17YoOHCCNZg9F9BePWTz2Rq3iU8oOB
EN94hEgVHTjwhGpbfowDkxJHr13BAoBzySXd7lKpD7J3PcbgtBZW+BmZZoe2MJ7fLoZE25pDkuDA
mMMpZ0Iqv2pqCIrsSUQOgyZNS6JWDjtbN8DlVRQMwmaadRNosPpouozek6YbHYy+i+kKEQUPnNJw
zSA5k80nzG9pCOWwzhh1nwq7EdwRgP3EGNwEZiIhIobvR9e++gCA2KRWMc5FxCTDyFqfWVd59kTy
XZboVUobjclZqrvhiJU93h74EPy5YNYLiRST1nfSQCL3f8A9vXyMhSf1kFE7QybJVGXjfZsODjZB
e9sHeVaESzwiKRNnsUSLIyuVMyvhC8NJ1mNNUSO3PNsnHbNIjGxEcIZn/nimqYkIiEce30dpYq/y
3jScbAgh2ygee3XuT1cbdDiW8gDav7U3UlB47fDCubrNU8HwqXAMnWELXHFRhseO2gEVJDu81MdY
kkm4tw0nckzeFU8yrCI/9/t1ikmjdZIIsJKMHBLqVU11X8c3+vYzwaCbCHIFcLLJOGLwLvB2M8Sq
xY4sFPHWHBpPqRNJq0Hddw841CXmqvWKM7VL2Mq+J7LrSQJ1Jx8ApdOVluGxr8TuKOUtVe5i6yRg
W/7zxaif4Lh8AQnTA0LY7/8NUEhF6iKpK8ahOlR3CoP5xiE4wgolm7LwwKhELCsLCus4T8Dd+Yve
Muwi9b1QaA4Jgv2gGXWFtSuI86LgRHReKpeL44ajDu7mfH7JA/9UeBgveqHZk7/+YCPGC3l48yPT
bsPle38IFuac+87UUrbk7R/pNqutbFxuXg5eZMpUpOUlVtenryBOSuuY0eRT+S8zKMxdupwHKmra
AHMxatLf5GCeKZRzdLf3WgVKZZDQ8GXQCwPvKOyujkyE2THbd2+siL2OHosieVyfN8yeXcCR7h9/
0eoVPUONWwQh2R+56/FstutQ0eh58i9F7yAZGVeiz1lnO+drkiHg7sE7MvPCmBi46Kj2Q/SOF220
eTojY+fbSgNgKgB+PA0hzR+aNh6A+vJCCLkDOFG6InrhPRsClxbt0yESZnkxZXTwQBB/i6LvEUHo
/ZKH7hEuTs1OY9/gHp87M/632zguPzpPx8ZQ1bp5xtB9fTknbml3376hPcZQNB+BU5/mD6KY9oBp
4/owe6qN2xreNsxwNIp6CW2jo6QkSFtGqpxtB0vlI0i780xRCGCDBh3nodhiScwm5+7qDfANeDNT
Tvv7X6Permqt4LBKA+iEFylrNldz/cd/sQvkCZH7QFSi3WmxgD69VnqNxIGtmqPDsSPaQ7Pi0WHW
RlK+ASOpp6ICwFW7c3MK1rFHzKAMX9wgjjj+oko6sldEkSh9mZHcevgboi+CcKjihTuqtUp2cXp7
dRXgXJPM8L8HgxhN/gRrYGExWYFwx3o26EClrCIdCtmvfABbzBjpd0fUim48YW63g4VEqm0shOVD
rcROHqee2kCyTnyx+VjfjI3F59IMoURZq/aUBnJ2m1JViZGSgcMGQnsJuutD6XSu7eqlmSeiGhNM
h0x1ge076nvnB2CgtZvoJu6zTVffZ6mlmB1h3A4+9K6qR6iFl7C4zNbp756boyoKG1yfcGlgjweY
6+igTbanYCN3bk/71N87WLuNUxMBv2RFpDfCoAtTFOQEPi5elcHrmnjCAOr851FtTkKagwLhnj7E
DBHJpR6z2DIu4reKPbFrXqFeywEsj363CE90VyWJGSpzpN3hgDqjjSPceC3Nbey7vtdV+b47nGs2
3ffd/1IdbCLlVSrZpSxG+AKwgKpitk/v952czt85UMHSdjwVjp1XdKQoL0hJW4OSEtJNQFnJpyVk
p9jJlrxPMv6VLANAar0CDR6eLTzR8nx762tnm8huZk50MdrTJTC6nPdBX3PqjAE1yIaVPK18ZX5F
uSBCRGR7YI6XetMQVfTZh+ebiebK9srXabZNfGhMLfP2j1MgabbhSpa3hVHplfSO0S/EUZqDA8tP
ExQOIDYRhLGOUUsrwPgJCN9hvNh0x0eZPDJ81L5e2KD1G08XtX9U73N4H2Ud6DsbXyAO5ySjCf8g
z52+eDP80Y+h2FisvI4DD7F4mxaTOtblng1OmAv6AzZq3Umo3WTYYpfwmuMe/McX5IGVmh6jIS+R
sztpk/n7WUXjipsXMl98ETRmfe0cRg1cp7Xi3rGediz67VGrMVmzKPy+ed9DkI7EPcqqNFrGM6DV
M63rAwTU2Vsx9U3ChpJirN+2XvcjYQ/DdiHYCc+E9fL3H6hW29yZuS3/IwM07eTJfDxqr6l5xAy9
L9qg1lZ+kmT2ktMlZ5RM8lQXdixE4FQ0b6PzmT5FT9vcyl/OdkulPvmX8YHvXLNrPpDwGLUU0nH5
lQVqgDTS/Iywi7J9MRxZ8/zpg49hOnCBK6dlDCJW0wCZ9ZVjrPXYZ1R0lytgPgrwDEQf0ibcVVhv
tCgK8aVGPFGe1HrJ43WPokzzGfLlQ0j3URjHUQVDYG7A1yjjQUAJYROH1fkj6fBKY0b8How0qG7G
bhzPaZpUWXKirZuIjJqtuClveAenI19WnijRB9yaVAGC/s1EkgCd93d7iXE5Psll5YyEd+YVp2wO
yddu441mouXHfu6whLLnMgTxgmOXWHvoBb5HC7VSSkwChiZ3q8lJsCma8VV46pwOxIo8kgal+JVn
MJOurFLv7NeWZx49XHM6CkFi22v2wwb6+RCLpVoLPuiHm+mtJ8DgoEWbWindoFgs/ouooI2B80qq
fVRxZY9yQbEKuSVHND+YL6L9AuxFIxyZeIq0sisZoW6hZtRLzCeB/UwNFj1P17tb3OGhlklzV5Oe
8VqAukZl7RlL9aqMFj7Jcwp3tMjiil1QCrAzxk/ahg6OoXB688da9FCXd6voEwCZWovjH046f26E
Y+0uV0w1exOBi1Q7HQJ3ruPNAh2vVhFlXj3v/Rlg0ufgNeaV/3CjYM6lsQAgDDa62ZSBhffFZVRA
cuS4xBp5ZWhx1kGhx/03iRdv/2HqV0oTd2YdH54F6eoBRIKBu0/WjYAIRVq18eqDydaGsuq8YdNM
0ZjDd42of/Kr4gneh2RTz+2Dwovjeo35nZ2Q4JB9ADIzGojQ6LzfKI4KHdXcR3d8cBxTpu7Zw68+
yMC6HA9H5UcKJTZPxim9ScXVrwTbDSOO/kwafxZ/T5Z1s9/phjxiz4ctBcEm9JQEPM0hdC9PXKq4
LEYwtvneYQBinn1cT0gxxyOWAHgiOoa2EHJEWwlakre3wZp+mRh0to8oiBVlpGldK/nARs4jyije
axyZOVUcNl22ngeMdRca9N7m0NIjnpfcjkDrdR+KHAV88jE0kNw4qgkRqDe6ZQOrJviudyhAFu1J
8ovuvlyDlEP0ITlCYEunjsDHludnCXK7qMaALRvdtpbsp8A1k+KphInB6+G+A5G+1+gspUcUz5N0
HuKU+bA2GMnycPWu59jmbfevzMqN7GIgMG+G6j89x2lONe1/MC1lnm1eZmwL/vOJyZn9C800AB4M
11d27pq7s1Ej8lwWe6rchTZ9tImGd2kgwGaXiUxWnc6cuODZW3uGzM1PShPJkY9ptAGPzTB77h3f
enY9DZxngT6xWVw7Fpbdxfa771YK34COnSFX1TE3tnv/yatfB+rX4sNuM/ru1plT0VKDpOrVhJ7s
TKboDFj4J+xWCIiPmvJ7/A5mVS/2TGSTucm870ZHvuiR6xN5Aj7/iMV2y+zF0/6yDrbyqKsihRhv
WZaKKLnJpg88T3Ny7cITyi0w3lYloDaK1LLnORzz0cJpvUIkPumDCU4Nf3YmbGLU9uP5z5/IM9Gp
jVJTofmeNzoDuf6AgXUrzDjnMlvrbLwlBZfDFAbb55E9K4L+yo1F3ez7h1lra+z+dz8nPQkaixpU
Lo/3sT8lbTyueDYtvFu27YyfJai7md3JxWkE9IYPz+YG1z2pe0yF0IIbgrRyPokdUpfP7eMkVk2R
HC6iKJRwQ+j1L3VMuXQOxaMMu9hQSBQGmK8gvHTIyUvJ41L/yI4PtCAhNKTTLGzL6q46JyNhuFnM
Oqdc4flAt/UZzq1JeBREU2n71DvjKZTfWFzV+YKnCQXf9YWyo9vDEBP+Xvucmy79ZwTmevLRC7Vb
cFE3Zzq4lr4VFRDvGn3CARdCMw5t6NpQ6CgaSOtMmP8a/HnDzeQYh/TJIm9xe5CsiQtNl2VGvC09
X6GK3UO7LlPOUL4yiVDzpw7gQoLH4xyS3V3RD6nBc6i8KaSD0wG17/liSg9kcU0kvzY4kj/Gjm9W
DUlFbEK3ZfbOyi4wFyUuyzS4T5pIPmoBHpnk5CYvazRTLkU4qft2BlD8Ed1XPhuGHbKXbdkZ6nDi
BQog/FS6kcK3J427O2aG4bREZ+5jVGX99Da5jpzbJne1Y3Z1ejQiq0ajYg5UZHKQK8rAJPIKJfG9
Rfmt+QD4nQpXUTyneXd74MOcpleRVccL+Y3/XQ8R+2MAyGXipBoYA7iGz9Rl+/iEeDGu87F4ib2p
+AU/DFya+VPGBdrqv5JPzpwV7Ev5bI7jbXqk/nid6syzAotJDAMwkXOWPlyXQdOjJcx/7kLAylXS
d+jTkZE1g8fWz4DuN4phi0rwvFUBDzP2ngFIumyEJZImJlFfqebffufzf03pvNTHmqsJc0efQImV
Bw1TTclI/FkGVVQ1jfm3nMSPHRnJ9VF1ZWdDvC7bCRDrHmazxHoO8fEHDDHyMgzHmBIcdWAI61iQ
Sff1Et3URS1+RG04OVDnFpOoALyDYbIaENZi2Bx9Xgro91L2nWQ33Q0S1+HP2nyOyFqpiAEhJdkI
xYFRqK2JraZezk3o/YfzBzzpsAX3HeSMwgUDtZd78M3B67mUBuiDVA2sq5AtmM3TdhMlh0lqxjiu
ooSjfMK24iA2jIU7VINA9mIjF0B2ir0DjxBUHWiw4vw5rldCHGDQU3WxTQU5pFL+88hgdva+HFow
tym8kTjwMqxfNHEFqwPdDF20/s2XTlbyqPUpRuwiLoS9NRw9uSFrqPU+b5BEIf9nkBKj3l8Md/3g
L//m3kJHXXCUmnRNZMbxs3EYPlO7CUWksCA35C1tDDKXqQ4L5naG0H+/FmSerGqUUOzuAtC1N1Wx
RuKN7bfH29N//DGL7ef1bdLPK/Xt8JjyvOJxvvcP8XHTOP7W3pbcUb0clNjAwQn1rOHowvNQhOBd
n6T2oWFV8iFZ/k1jNorVDAiEDlwgbGrYBlQMMzmBRd1JTKb1Undq6qUzQAzcIh6WiBbe5oBM0Ke1
+LsgyKjkgxsntIMUNJYTfjQg3gIhxillQIKoeB/e16BS5Z63gPRPT0kGwAb5SkcwxDIyLzNultJE
impIOcUXLCCgiNjFlQs/23oZTRttpBh8x4dEuQz715UN1JrSD13+HdO2PQmCzskteEP/Wj97Hhe4
wRgenY9tBVVpLE47S2ZPlm2YmTJaTL7zIyPGZZUlAfi0RVgA7klW77l+mCdaAc9RUy3KhEqzMcLk
/9mOYBCL3AexIbTootslqFctoAhgIrdQiIF3F1OP/NE8/l0kfQoqZvdIVQhlNSGpC64lZ6oBhSCQ
SN2V8XLspzL8dc7lTI+Ug17wmXH7QJoPXA/PRSgaBsLtivGmVaLzKOyM2OJnG1RE44efNJozF0iu
qYMYm2LdFKpXBK7F15R6rrbaUy6WTNaKgp5lUhTfr+vO7X9zl6hpu/96AwXQhIWL9RWKgpkZ9PCC
SJop831kUiHpH+WCWf40tUW7uEKumOCxC+giYDQFA7elB5vTYnuPyokQkyPxQJw2KcGZpTtauNJ+
djSOiAO2fymdRJ5tJl+Kw3561QXLEjGLpn7jP5VHYN8UH1o8VwUXaXXyDMvWGBAZeJj+Z6vTq34s
RzehFHOjVvib8jtEY7vH9pBpzV4pxXnWvb/67MYHRN6pdp5LQY8CivdQebgvT1glnNqRPJuzfWGT
i8HfPnBuTyDvfRI92sDlVKUGb9ncxYzk48qlGbkXBuSCn/BR+dQwUsqW7HpBl9MhO2R69XQ69hTC
xeClmRluYjXJNAGcCq7pPGaJAz6Jzbv2xAxussfLOcnSx+Ho3JoFYQ1PVzbdT4echDdrLjfggqUy
40GGCIw7Vnm8gZK2/i1TG8xpu1PXuwo+IrwCu/s6NGGdQ8DhbUlmInE5yxd8/f18Gpm7v0vDcQdF
naBlNgLoAo20xLFWizGmwVRAkgjXCG0g67+svGC+M1FmeAjiOEMBTBu/CZkceC7iJdd0yQNup4BH
BQJxRNJK9AeGCRruTlZl1obn9cYkKYWUyuR+jip2lwrOS2Rw8QX2tSyU8ybK+Fovz2glS2rjZ+pc
FjAhDdZHoLKNesBkngjiIuqkfsQHqFvrDBbsMDjxGG8DYcONA6GiAA+1VqqSCgKX1PHdBYIhUbCS
VsRbnlm0SJcqK1M1cjqgv4nhohfC9cwxlZ8cefEkgu2q50A1mfQlHUwU2cVVobxuMZhW8gkuejck
ZMddbk5snBzBjVa1IgFNguk/1sAAtPqoZATTIcJTkW3Hz400XT4iZfpBac+Nlg750K/UkqoDWS5B
F2PBTH8SQjEdLdTdxgIIGV4aQu3XoynZoTn8Jvz4IOSQNCiGPf74YoUnsnpkp39+091ZwSWCPqsY
hWMb088tnXY96odF5W77APg6q2fjk6y2m437C0mC2B6ssL1/ZOfC735/POIlcGvRFIg5kMzxGsE6
9zbDA421RJI9CJ4knLRXacmsN/QjLes2mK43070+wb/fjDjdowI9Au/KG51gthdfVglAXFSBvg8f
aLp4RJ/AR+1STQy6N7NbtevvenWKKWdT4O1S39vphJuvD+hi2WNM/l1fzUuaC1NlKnfB1X3MACs8
gGeV/1k+YejdcADkc+U4NkhfBQnZJzIoIIt9Z1F+q2rZpFZs5OQUzAOyG2RMWu0a/BzANU3ZAfkB
aOwlQWY17CAMJiu76S73jfwF9Wi+SFUfxoKHIKbcwRfdlbuLlnrhxQXE+dezulPK2wqv4bj8yH6Q
Nu60d1PKGGblaZClBcYySXJsYraX5BO51dbMv+lmv7bKfbXkDlNgIO1uf1MOHoLEPwR51L9PSlwQ
/LJvwUygom1bEGLD+aT8tQrnkvSW1IAXVygRFWJbYZmn3QpdU7zEYxQ5u1MVMRl7BW8v9jNM9jZI
QFMRAZGJJPhNYjEQBzLu814ajqN9/1ePQ222x8Qp2zZIw2njD9+vIBGN6WfQES3zJWx2US7wEBtr
7Bk6GE2Q2pLwxdRBiyaTcwIaV+s1paQdWTRfYWqBPXdXBZn8zPzc/CD+67k5VEPv+ZwfMAXW3mHU
mJWKZ5zcmBovKAKTdfn0Q8/o4fPIdc1Rwb76zBZyxoA2pBeBMTblFdHHIZTgeGftsiNYVjWrNEwU
6e9Azc6J5XmKONv1aMCD8u9Tqizye5IU8vV+W15Drd5zVWs1EI8jlmgS1/5Iibex+FpD+qn39JRE
QwulmSDBa0YEEC3Vm8U0ahYQngprzyaXN3hZzF9CedxXnBXfxLgoYH9XRx5S30e4V75C4DhVD58J
BuL0BOVFy/WnpTzJcgY7JeSXhf+4dcM/9UzH4I4Ik52b8sXlyDxYw1ApSEBfDedNu/zgC6kkXRaj
z2mVJm+lDrdiVxmprUSgJCt0T3fjujr2VdEM57SWiV80dUCKLuoPvU1r9Fir44Om+aM58hoID7tQ
mL6Dl2Gg26vQJLlnKxO1ItR5Rvl0+jchqljlOJrwKc0fniUOPECTcybhMbZkWiWhr1MDfnhPTf8S
V2uzMhYE7Cnu/FGGzWoq94EdOXlstlBwTRlzRQxT5utxyU1yCYtjnre/R7jF69knQLdcqDroQt69
W6MY217hg9qUatWxj8MfF0R0n9g0KzmgJCZ2oG33JsSZyoh2nWXYmgT/y58f3UwitWrb1kbRXDnQ
OPiBfo94dg1mwbr07nUO92R/UuFHYAcSTgoimkxdkmV/rZAuzVo0uybtp/++WY61oriNv9Fq4o5H
neCkNH7iIR9OmqYkR7JoTiT6SyCkLtUA20f8ViA6ix1nlU7uZDyqfPMnBqzD/R7JpKuKjD+gKFyg
hIEEGngMgptKplK9ynALVDVW8hzIuuPgthCSbVysK5U9VNU7QwZRcnyvamnPAClU24Al3hzq6cg9
BYsBB+Js85VtP+xdqPnByEQ8LhUjM/6lOvhZlCeNOz4zke/ayZpDGiS0zMKw9hUsc82nMO4odM2X
hPSy/UyQIUymxvtJdoe3j/HLX7hrBClwtfbvfPpf/3utmIvRZBSu4D1OniypfdMIJUCVSZWsjOoO
y/NslmkIqDMCLLobTfOoRqG9D7+Q7X2ondFkO+BRY4O4FiW5Vq3oAOkEsvkYlD6xbT6BJzsVT17F
o472fSq3LMzVTKD2j6U3qszXpenc+qfux0MzGWownV+gqTLlbRrROaSU7MJ+MSN9zzX2n4jXVS7X
ydUB31FsmTCU/ciH9fnGWn3fhggypn7a/k4D0yFSqow4UftHrdpJX8XzIO2b3CoE+o2SZ+v+pSiw
TQ4sB258mhwyZSfg+IM6j2h4AXm1ldgSUian6irqoH/EIRMMJQhF2tFjGXiSvDMWm6h4NiqkjZ3g
lE5vZTmcp0CShf+Y/AZjUYsfY7FdKhU6VD6FWxKx/sYgNrC1WbspTJFCazoBWnJHvqIzF6TswMiT
uMPktazRUYppLsPaByBsv+w7SPk1b3+c/5JLECxV/uO7Rg6Xp++HL3rpMPzB/06jcTOoqKNpKsyj
GHhdHrT9gfi+MbhHOZQM6nBZB1nIrmwIoeGFgg/f/AERHOPKEqlj24tsYYI24m497DJvVa0JiOSO
retB71MRh3Kp/mXbcxgCvDew24ECeYw1o7lp/7ym/LyBxEpYT22jMDB67ReZv0AbffcgUl1581zq
H/aaXr/GBu+JyCRVrRbRfDi4PY6TbIvX6bb1W+fTMIocHM7htwR4EuzS78bWH0KFrrCDBzxZlH8r
Ycne+1RPP5iIX3v+Uy2+QM47AfXGbDzA0oX8AKU7h1l7eMpccaKNRyBwr6IncTEwPxNJz9WndSds
WAOv4UxSkLTk8eWZxNe5eLLavrSIsZc1W74IZUHjRETBNcYBcYiPyc3l/ySwHjKxG8I0jxgpHYnD
eaG5CxI2mJnpGWvtwPr0K7skB8LE4fpdJT3z76ICsoDfe4XHW0X5UT2ldIELv3zR0lnrycLdQkEO
nhzAy7FYT7yFCyOgvg+SFNmdbBHVzczX7JUNSvwEeP8iMyPIEFEc97TLbleBsjpbuztGjRjtyYCl
tuEmQ308bNpi0k9a/K0y/zO63aYhJuJfAlUim1g++xIZ6YCFScmKc5O/KXK3ZjDvCjCq8Y+cQlhx
/cy3tT8iR6lbrt5PYROVXOQx4XFg7wNJUerqFGeRhTI3tqyxThWj7spE6ZiySVDdgp+ZWxKINZoG
lROb/CP27WNAwiflkaCPH+AAwek1FqybLmK/1Gn3pUcl4x5efTeYrd9vQPd3JAQ695KxaCNyXKKs
jAQsLyAMbPExYbuPpZuNHGGOQ7kVAf2xN0O+jcqN8Fi7fr/t24hoAgtayy6ynj1hMDOK/plbtzSZ
L2xsW1WekeLtiPNb8r5tpVMAE5kZzoTGfH+pyoLluE0+04FI/0t8BguZBe8U+DOzXIIg3urStN+j
CLD9QOJoxJDGn/NybMTL5r2c9ClDxabdpA6lNuUaa0oS5KEjqyth4n80YNqfUrS4xan8wFf/zejT
3XGZDhIdvHL5ErWfp3xSTMBjdXtKkxs99I458YCJ0r36pYUAO6wOJ0djDYLPBCIDetEq7PF3iuD/
7jS04SKOskjmmg53040ApOfbtlgV/ufkFW09Fn+SdLOm4TT4avHT607EWBQpzGZci+adBZ7riL4Z
x3aSiGJxKS1SJKvhiIAtbhJ7GFY53QSqgLSM3MmC7vS1kwu7/ktlhHDGRbDSnOQM4JueFWg2+FmY
PpBdpWxGRzHPCvKg1jx1HRctgc6DrthNYd0F/H8joItme+I6GVT2JfyrJuTy7HnJHev+id3KNHJQ
vRquFo0yAGp3vuJhuLzlxC+dwHW0+IyyljQ1dGIByitz0MVeKz+n9perJAd6ccx2BDai7QvQwSE8
dq/zhh7eL5E/bG0xskPkBa/+DAmqVGpv4X/MXFqc5e5parFzm4IqEe5Qh9zX5RvgWrRkDQC3rtC0
gK6+faneCYTNlbvyX+IUsbF4wLMWEd+AQ7ROPfSKE9N0AdM3ExLSvU/1Etg8DakTNc1/8OGJ1Uxb
RxAXe7r8fl9Dgo1t2AearmAKlT6/j/fUpV6It82DHhzGJ5j5Pru57XdN/Qp+GMkJ4yosqFddIWnd
EyEXgc75LFetnIX9qkW040W7Lcxu3KRazApAimiVAuP2pSVkKuuRSnjSlaM1dh53NepEldAqyK69
yGBJcGrQX2vsRCFr6Zt70/s6Q7E7LTRBNGINTZ49+u0XzOh7AfWUEenMAi1ES1SUIbAmCjfSGgD1
/k1RlK7OkOPBGOX/II2xgQxOThx9uvTwBpXxOmtFr1G1YoLrazhHP89U++IKlwajXfPL+G3K7bMr
X7MQIS1MhRz7x56qZ+zYgr3JrkaH/OnedZHblfXQ1PIuCoMNDzQ6F7kMRfRiz3DutSFOptFms1ir
qgg8KVDr1wejLQFhlNJXsfyTpzZJbrc5rqP6Q/mOrSNYxEPVO7DBDMVRlSVNfKTdqG0urvXR4e0V
zn7I/ZBZh2rGxHQjqAMjIaCzAhL1A42CNJcR+620K6r9LpC3o21jLefyS7EUJuav49EKVMWT5oGm
CIoAQ/6nM0bavPQENjE7auTNRH68OSxLpaP7/vBZV64ZkWZZ7IM9L8OW2d7VS7RAeiOXAKVPvnOh
0yxSnkE5sQOq8+1upAnc1OuWbpNsD0hgJtn13Mm8l0ZfGkcEoU1xKvz2gNyiIucTEybqiDHQDLvO
VKuE9FmhTAuHaN6l9GHKf5YZ/kzQ9CjbQjRXOYEf+mB/09mRJ0LKiEmGboTVFER/KOmjZ7TqaeCe
w66zoSAcooQ9LrcvLPGYPywCiljTUkQhx9fVrtyEnVVHsiC3CPidzqdlNkMjuDBYqEpDoKBqlRmy
zGo6hS/jDg8zdPlaCZ1zTQYfb1xQJVvuPSaZM24sN2NrV/p/LfjQd54TDXynNqVnJSo3nzQu3MOA
jqY5To8d49QIh0jRvs6xMwV/dHuyuNpjBtBSSXSabmBjjiyxYXKVxKUK/UtUFU/dYfveWFO5H27k
6UXxRVzWH7lnILDLHo04tq6Nn+3+bknUkpW7RwiRmOytpGZ1BvFT1PbDoQ1GZQUOMQ+keMkpwuc+
Rs8q6Z4u62y8s4CDssQt30tWtCfffIhEr13U7LQGXUrdnZvv5DJz7xpF/n4ulT/RcR802F5a9PFj
6re9t0h247HRDTFFgR4qkbJIiSyI8CoQoFluuOF1B7UsqzW5rbLSZKIoy8P0EW6uBQMfrqSSpshl
QVX/7lNRGcDkMNhzXivSJzqOKg02I05pMAJ4wOcIdPGPQ+tKQ24aFHkWT8yz4AUzSdKXKlm3Tquc
I40x1xCNgDkvn6UWeoKD/KrTZcXeBkXLqCx/UWQQgbJ02NSDvutk4qzYjqO9MImbKPxvPchXHul+
nu3tyjlrbul0xpHCj5e2daq5/8RTWeHKxuyAyuOUvp3WWJL8KKNc0Ql2K1pkl0E+XbVkLZFIxP3z
5tANO4qFqoNHOL8maLz4bliotGOHxRuV5mnZLkM9tJFsQI/fWvBA+SE95Dutsqvmcs9HD8bdLGP2
WjICUTFcQE12vW/mUCxxTzaeAfmC3tTciwjDdE/6ptyzJhA7R5yaT9/MBveZPPY5A6wDDpjhbrgl
vSYLZxNs+4g7r9+tDjb/PwhYgTpPED7vocM7snYjVF0w6rIFkpVrzVqMjHJBts11tZtapAW0ri6B
9F0q6GhxJjDMPAznmFsvyXdLV5Js2pJwANnJ9M7hFecogzhP2qjF1eJnqX6ReYBRzs/Gh6l0zfA6
ku9Ii9NESY8hCLHgzAoRTPyUkEJ7Psj/rGEd70TqSIAnmmwlzlrcZKgpT5wIYh+WNIFN7A5ViHBC
diRC2DqxyXjBEkbHRSuBQGS2IWrX8Mx/pj2IAwgQwZ+oyW+f+vMpJRN0SypCD5/Ldf71HkoVZPTp
gRiOmn1iwC0HkDdXBVnsSb4o7zH8GWDC7y6P9xiistClBmYbgt0b2RV/lIsQ+Ad8AzrPbpyNlgHk
ud5WE9tEc/eZsMDugnF110P+7CdRA9rw8xHeLZ+bG47KTFaGQ1F6z488NT5NU3qmwRKHUBLbHF4O
jlvKuMOhGITrxAOcSvReRhXchxRyvZbnMUONL4V3xFA3zo4KT3iYTS+T9Gu4+BP3AeoAxLjJPTqq
fMYK9UC/KeaLOle1W2DEDH7/M2eExYhrUTDoC3OosDfUn89tFNDZyr58ebXc3Y4HKQq3hP2y/ai4
GrwzAAF9DFJ+K9xUWUarGG6upZyGg46idxVQtsZd3xnzx8aP1zrozpqjbipubCmDf2egICGNzfd2
y3NU03PcZGWmYFGHImOwzin+XAfbWl0W7sP4axs9s1Cxrb/z2CWw4EkTY2xUvtA65NweEMD+2qKB
pTKl8CToXeCi7KdnpXOO3m3Xgu7l+aihZk1P5+vdev7BjAoQnSlAe8P82rqPaGh1okUaRDXWpSnF
9Qv91W2BLkjEVWf8PHmilvEsKW8H1Yp26Eq7QAnhPBSSii5sy13gS+qhkw1jPmElmx/MNVw+bWbd
j0S54Qwe2qO9Qby7Fi0c8+Yjade1FGQFkWZwziyFMW+Sqevo8oUAJ9B8nCsicWGXoMqJNtBhtTrk
UdHatNYVa4jc8PYtqMld+FvgFgjuvy4XJm2mSMrAWZbWw+yEI75T1RAy1r7u2R10FGGpUfTXMhn8
rNHa24qJb0MkOekW8EvYpj4Ru5ahjqNzw6AjNoHV+9OrjeH3FZGBHEK/6UmHTgoHLIHJ2QlMnpEk
+vLQJ3phYTqMm+rnLvqnXgBjy/NDZpE9uY0Taxk1Jh6PKjTqGntJsA9aWzKNExFD7KSh64jzJxVl
OLWJvYOV3dz7cUA++VVlPjaBP2K9Du6P/S7EVbKBHWQ2s7TEHPEaBwAFLFTsNecwkANcNmATl6DY
GYfxD48F5R+XE6G++pxOqjtIUTGFLGKTAegmnFe9yP5tT9cEQodj9rcWd+OZfr7aabwi2NIRvgEu
9lNzeu8RWti8+cQNHS6G5KZsLcpYUVE6W4UJz+JmUcvbjWrrBvccsDGLkEnWnPV76KVLWtTLZprK
d0uTmnSyDjtEw4TZiyb51Db41EElH7TG2yWBMz5T/MUHDHDX17BQRv9mfpCsPSnxzS7p9NylProk
x0kQPjPDIBqnVV9Rx2lsLXy8eRMXIzC3JtJz9iz+imvVsBS1u70QCJWfupkgAnrZLqIh6WKNuMp3
iwlU9BGbWMud3CbcnzFMIQ+hxIJKWkEE5q74QFxoFXh/1q5JPnSYo0HPboPN66H2V12WkUTlvtKs
rUdeopZo/t+mKZlbOm+rmVZtdNks/KIq6WzN26VpOS2KMlXwNsH6Y8z3oSVizzn09NbH3okebCDL
m0tPjpVkNv1/q+4emKHgnnq4B5ioH9eqRcrY4XxZiPclSOf7RT0DoEg80n93kpCFqhjpT5sdAfw8
ZTf3UiuJilrDX/PxXQWtsiR+OHS5p7Qwn6DOK1rtIlHStc51LwFhdRh1YIwVj8o5YXsBgVRP+Eni
8LvclCrMjbs2nh+2aguYD1PXRSDQWMzuu88EFB9Gfo8acSlwHhk1J8uPvhFnjn4+QvKDUDYqlVxJ
7IMTEGbTIJpS8uBS51mrU+YJOOKtYXCbztqsKY2IldTL7E1N2Z5S6hTdJIr3oVc3Tt3ci0nM75ww
40vQl8BnC8lI3l5W1izIbdvQd/Go1jblDIxAliHvH0AWynGv2FQl6HtYFAxyDbQbd5bOeUENmpLc
KN90OKzVAVi1+pWYnZDFcznmVO16s7OZHmULhUccs+lKI/FtdCmOwZC06IQzjI6qoDhvF+3IVn8M
fDf+sTF5sVBhwnN0GaDnogf+KEsMWTpDOaHN8Kxf7RmvB0tfT8N9UMHw+l37IRica3oRwZKsnjk2
pfANHR0H1GNuBbDmaD4TUJm5LeHAcXxC4SMS597HvlG1ebXI6KbBhLD1v7IWSwRfV+VBguGKOdl7
vseFgcplIwVzhUm12NyyH/t37bkx2ocT4nPEzQ77dxR0u0uuv0d3H6DAKN4nQaDuMb5UZ0BZh8Ef
Cg6GNnOFTeXV7weUI+LN0sncbGx09woD2vYpoCOkLlIG1WNGZ6xwKFXPlAwZVeqCin7Udz8YRkmZ
Eks3p6AiPdkZQ34cvm+JtdpCP2xyq2Fuv1JKFinRdIHgwOVEEm4TJWF6Yg9aZqtRquPdkLyqDpqZ
r/fToxWmQTHH6McvNNZ0C04cTcH+TEOQgcHdtIRpSRODXujra8DuyJucxLoEEmf8HSvPJI7MVwgp
jjKaeHaXhHVsuh+g9nJdcZw9S8satC1MT9bRiY5mgSBEf0WaPh2+zLUDLap2wxRVkXM1fDGiK1gi
RkQr9Bg238PFJ02W9f2pFrkO6BnxV0V0xF0lfDpnVcM9Ev2eRkugPQOsJjseFKTC9LPVn5EcFqzm
zMNhHI/hwivhP2MTxHRzTX2i2ZFkpEVstxDmzCj0Q0DbYW2jk+lzwgmAFMbvOny8HDSZLUFg/KCe
Q/4KmXE3KuAdsUg/r2Zn7Ly1Wgd/TPunZrEOAHP+LH1j93UDWL/UC79YAW/HZtsdVgyFI5IpuiYh
7EAuk5nqFlbzcDUqUZY+D3mZVMy8PLXe7Z1ZKtA1t4X+xzpLT+aMNwtkSJe1HgMMNZkHKHQzejcV
BRpOKsBI1YyoyGRiS+VdGqIs9/ud3oN/CbXQk5KCtVDjxqwyQJQ9TMng9edzEgxK7dkxDkFX0TAO
Yhbx1udF/KWkJMT3CrwWem98loKTJI0fD3UEF6V8ig9tYHwjxj9gUkqvL53ViS1CPuD2bPDYIi5t
DeP6ACLPg3LcUatpKWyFpdWSRMHP2besG8O/XMgsF0zezEgCtKS3xqsZJXDsunEJh0MKASvkFtRe
/aAv+ri1zlP1PDOX04PsreHYjfB+0BktCSxrtPXPVJrhRTm6WzLmbTw9pmWPuG3OMqQCa06cLifn
91m0KuTCU+4vYIlxeroH35SYKCbUouww/RdOBbnDA23o233gRg5R6JUAwfnLPLtObvyLaogMzM0t
MIAw8iwM7Mra/zpmKNSVF0A1oreicwobRfi314VustyLWWSUM3OSHRl/TlpKFIo8lPsajP0tMt/k
7acHBEsBrfhvx1Dy6WXLXVh0VERedE5tXeFbwkXnHew7Hwx8q4dLjYSgW9tPPhpu6in8JNke9fKp
U9iUglcvojfd2qV/dw5mQlEMQdDiK3oJfGK+RAjbxQNJnvGYkTZe4DNJKu0E1+i3DvgY7th29uS1
xvRl0rl2jc0FEqbhcoJmxlRWdTRIQnsTfdG97U46hFjBLSfzxTVCuR6mdpfMgQCPcva7vyU6OPCY
XWAsDTCVmuV179lQCg4zgQlVFRFTWJvpa8ngW9JfIy1bJPS4zinyCDQmrKQv30shpWRjnDBWzLnR
QmL8grWdsmZ7l39OD9rUMicmvnsCR+z73ANUQlSESsgnWP8ZV5P9V6fT64o7FRKvLTFxAHthZVqS
NMK4VUnzXjLH+xfuQivDH/8IUEB5WZd87jbRInCdPZ914CTsiND/45MD2Sna71ZnBiVgfuv/Ok2Y
2Lhm3wuCssyQId4tcqRqJE0lrQfHngQXKjeEGIP0EVEXRUve+7sxOnset6Sb9+NUE8FPh63JvNzb
7BSxSgI3ullUemQ6kwjxHU87q8rulykHZdxbQVjjAoMk+Dwep5XFWWmBK0Z2a91wdczgGkArGHJB
W2DhYDknNjwb98Vibjd1i0c+8YASs9XsIxirccMryM9+1awvo2BrDGlrR7Anyyir/XSpq82XGTyE
OfYSOE7fecgaWvraypYXuJDW70yvtP8azZ/asLc/ngHIyl64SGUsnouPu0Uedy4arD/+lk2L7SDk
5NNN+NrGSZdBchHjKKLFtM7IARZ4pyFxerq8fQwoSXl70nbKMd6cYK5795BwLXkOAXBCk4+Xt/Aj
iOjzVXn0fBmAMdVdWFUNU0gTgm3vgAog+UHPX85GOpYJeqKkYfPkIaJ8bAF2uQrDoDiPyUzbUci7
vcBOIK0OAhkcvIuTLDpmI9o+LSMsXJfXhUU8biCxfnxR62UBsnyB2Xa20N5u6gGpZcvo/dhAOMD5
pUW6gVUR1mfL/W4H5D0uMi9NeAwSOSLNezaX++cNDfhg0vnf4SivHPJHLk4URZXl8m39OTALNWlX
o2pvUvlAD9lucrvXj7+Wr/mr6+1gSCjDdwXN7ewJwwsXgkXQsHtawqFW0UJfWL4TdUS91zF24ryo
7sKsrnd+vFQfoTrwEE9tnALgKTFfFSNygV5SIq7zIQAkbeNPXSFrI++TPfWnrxMLFNKc2oG5IhL/
d7WagKYzCHKaLQxnXxPUYSVb0BHLz7DQVKYoFnY0XFwhn3aBNppuBN2b4we68itZPnRFtgfVI62v
paGUVhqzP+tgycuj/U22/n4T7JvlmFUXldrbuVAB1gNVmO9Jla6Zxfa92IwFTN27N+SehVG82iJy
x3x5K4czk7gIDiyqcHksS6DbvtXWRE9tEFEr2vUJWUt/UXwhV/YECGofd+Juw43do0z14QqXz9NI
UeXWq0tmwCw5LhJ2jNaDyatYm8n7jqg+hcQsUapf/2ZUctshk8loEElIart9CQ8UxnG67SC/roq6
toLC9oE01ElgEz2i3v2iQsVFH3Kn4wsbIJV5wTY3EnSpZhfT8BVslc9Yo34URzya8Ne8tJcxhhJI
gWO9YyppGmIoWIHJL9iPKKOVkH+oBNoe0W1SS/R85XKEnL9kfGROp3BtHFEH6b/5WBg4IV6ZyxqY
uYQrSKCaKzhiD16q0nU/h5tGR1xzXtRyWAXGqLXUFx6bLLPdIO2i76Uhvp1tIm2XB6U1x0Z+wSll
K+A8tpuIyiM4GxVk3AXFzQL2QXk89CoboPdbDRvSEcM+1LSeszgdFVTmbE+8Cep0zcWW4RelfB+K
rDn2BraTl7s5rMXSZGUW57dCBagJtUm2FQmTuyMJiAF2Fhvq+5PpV9LuGxxmgfnmnLNSMmVLcBLr
lpPU9O3t2eXp82bncsMVf1sUUOqc8kGscoXIhBqrwTSgspeNUhRvmKdpTkCW6D5SDjtue+BgNwMu
YFFLYiPyORYklJYTj2QeLtSemz7399+43zM6tOCA+w70jhaa295x+aeyvXzvWU1gu5gfnkhlDqS7
o1O4p6qHDxYjNLqoEl71SsC4KbBjlydpekBPCYOZsnzfEBV4eIy0eQd/435sxKVRq0Rb+oL3ZUHS
z9fOHdIOODsx0YGyaFUNc+bP+z+PP27anhbbtfCLuiZKPuVG/LWoMSrVryMssj/urrWV3fLPSWpf
MmTMhrQTUzzmDQjepwi2NzAtDb7K6WFON3d5jQN09TOEiph7XlSPODg2ZAOO17PIEe32AI3+38vB
pygAu5C/oORkfeYwmY1iAD7WO5Y4braWZoBPu0eETP6cuMI1VjMCwW6gJTHvYzShBPPsBghsBhwH
cQyb9CAxbw9VztFzCRMRg81uXiCb1WeECu270L75yFcFozsITtCcpL1BFx/WzAboaFxm3a4eWfJc
gPYRuzXuyQy9SjvDoVcWcU3KdLmXDaFLOJU1EpbtdZtIMnEUP0Sa7waqeXVg0JsS6aORZX1iP5ZM
bcDUTlg3YeRuZcMAiDT9fMaE9GkuPXhTN1f5QtvieiHKH8cKNHbcuPl66pyKmYCrmQ4Hh0jFFxs9
OHNMCmzV0J9cqH/Al9HIluBN67f2a04HBCCrCuZt7LzR/oNTbgbCKImZ3dgxbSqZgBesRw/IUxtj
XgCW6pK3AtZqMaalwDJxX5A4ne8Zo+5CjqSzpq2gX/FUL9WrG750gsbdzwut2/nqLQPxqz55yXUs
eLerp/+t4RwFr64BUG+dfxA/+Zvd7D5N7tlf4LBOv9UApTjwyxFDNsYdVkIy6hI3s+FchsYn/nHh
fTz1rtXbU+PiP1QQY1LYLQvuW5C3NhK2eUTpq9Bimp/LdgoSD87oPj20vNK4C3mMjq9n4EaBbH2w
4akZqyc52oIvEaKBobbhvWLijY9i4VBGmz9WiyjDtzULz28uqMcw2DfljEgydvOCdJTa6k8q2qhs
ooboEwj7I3yQLs5M6ET0lbqqiOdD0W26rGFTdh/CTQGudbTCL5WvGcNtcZGglW2vj8fzDxMaKfcL
/bJ/TiMO07JtcRiMgy12E/kWGRRJgbPROSDttBG/Ib9l+CCkIawU+7v3XWHHg3b/RTQRbaEnEA2z
qONuacGediMudZqfk8SY7VnjsjST5LdOSiUBjAARuUN6x6m77XgkVJ7oRQusq3kUaLIJHpSnxC+V
BgmUoN5CX8qnF6gkmqu9Qj64vqtyT7s0pfCM3wdWoPKuNkCvMxPqzHsMSUgtQAgYF3AXqOcL9BHe
7G2WPWoZX+ReJS+YV+Stop1CKo7VCJFx2hwFDd5PchRioLRX6+l7roOy5UsUBFNW3UTczrwXt3jW
HCAsWDDp/djiJ1wPujvIJNpNPB0UPAE7f7/exiycFIWLeGgtIio/duc5JJpbM1H7QUaWapF8SDAk
OjxozqhiXTu+mevcRi1jdUf3Vjb46WzM+X1eTJ07dI+4Kzl9ey642yAsArRF+oja20TfR6c0rBF7
mBVjZ5Mm0ew9HYmwMz/FJdnH8Gmxiynhhd98Zh/ZYV3QXBMhheXW7Etboq3tjHfWPkVdvrhuXUHF
6ZYo4U0X7n46SusP8uwCLieGrw5Coku1FM6QVguWDTYRN1c56u9lZOkkmc7NBCshmPIOVFtIAify
RpG9JSttP7nMvmDYr+RBNCp4131vwwl+uM3p0UvtJWtv+KE/pFp0FeaV5SbcSntcmlN9JJEWYq20
IyPxEDDfQEsQWUprj/fVRnxiqrfz+pHZDidJKs8ZC86EetwDIG1TxfphiXDEtRKpP3GnAAHPSLN9
fMSl4J8w/qGvMKXeCFE1+838K25EchP8YoOHUDCQAreYaS4vfBOAoLHb7AxdHwgDibh3AcdEPtvm
3RQdTr0fPF/ov/lOJVa9reP/4lg89BR86hvgY+8V+Rm/42vuV1I5BjqVXOtcE5Xbu9WQc3BWu+xW
t4sp4zMPdscinMDZq+PYqGE9Noa/1VsK+vRbUnctDN6DSSfAQuAQlFu3WvXIQcAykpfCbK0meQxv
vtLazVM3uk1FvT/seMqzRUGjAw34BP2WLkG4l/jUuWzZWc+9ba9rlRW4dIcbBCsA/OdGue5XfClC
iAGufOodzFJSn1Qu6RMRpSNnwZmxbZhBEAglG2axERMFWSXA3OT44fU66P3TDXke0yk/8VKDYNaF
6NHLaF2LaDeCHQcsT+gUrumPckJaOw96f7yUOchjz9R/tTT/gH1qCyZcop8IUzqKXAm+2ntcrpat
jlONtmOZL+ukjdPV8S+JE6KMyHmJttpu6C9tBWTHPY9viM/UBWPipJQVmQZYuzjHG3YBraWCsZBS
Ricwlim0G2NlPsgftFd7x150fDXEQQcyDV/dafIATT1zPGqA00cqtAT3W638S3NDehtXsbvdXGoo
ke07qeg9a4Mw8zAaGKxHLfpb1cNlUixrelybSHPTiRZKaH+YWqSh42sSp66Z1dNNhS/6nWL0sIAm
A3ED+J5rhZq1iCf9wGt1+23kuYclphjRJAWykjTsCEHtGywvfdSd4i7HVQj+FjUJCjSFj/qa93KX
mKFv5b5oirkX+IGDEX0Vi+pwYwIPtm4Fl9s816CbDOXvmqEF9l9ekhYvAeDwl9/JdZJiHN7U4DhD
5bhWuFhIronl2AVl4u4r5Ene/tzvXWLBAPqcluYh+OanmBC4uMHPPVmteQGYUDVjeLwCm49zjMSC
THVyoNhccMgvwi1zcr/hxdBYN71LNzfFbSYrJr5YZKKFmp/eWnL8jKAyPFnz993AkrA8MPYptm7U
vATykBfE+MnyJR6iJsKNSQpcaoabzn4TQOqGIMM2W0IEmcMnC53Nhu8pK55rI4yfZOgzVeg80TSY
QdjauxugSku7gnkrh+cbhl4flJhJkcoh4/tkfyfMkY5URqx5isdxnXVnlqldIoy0OSVJiBh1E/nd
aaQCnZ8fPTZTdwYFUFF5twCO+nLKtTFgRBjU2tRpZ5AuXnWjoR7P20O7EhI2vb3IF9b07XlLpRe+
K8DpcjI3x0Sttj2T1E8rdtB5YMzPOxL1RnHaiKJ6DnzwY0sy4PD1gmsCNKw4sejlFiML8NHpRRNU
333kXApJCWPHmvjcXLOVP62vQTPeCmhODPrkTnOhOW4zXBqSAA0WHluJDadi759x7rzlfEfk24Dk
axR4U/63084lA9NcmoSxL+teXAkQhQVLizW4zoUl0DvKmiR0NHwHbhlNlTp1h44zagiEJ6IunndV
LFrm0/uHY1WcwU5JnaLRKyRBReipQilukQkpr+mjujmGxzrhEiW25LPUB+9tznvIwZ73F4TkyS/H
/GahLVciGaGQTpl2gaQTqVGDlrDxZ1uCD10x1CdN1LpW8c3qP2cI6mzwYvFoVceQDnVLBMXmvk1x
GDmPboeYzvKCOut0HBkFSbf20ijS5btUkfD3ig9AVaAYTkpxok6g4tlTHno75JUhh6RqnFuTbegF
e2bxcDLeD+najXVjEWTyYm+MpqmSbmOLHthsS3O3IrDXnDdVUAYGCvdUsKo3ofyujGdVjGawiWdG
SJKgXW8Nb8sCGaNnFp6wm4n1PCm2GQjyI8lIP1VKlkJkj44P712AYpqBTCdxyOkxxUCj2Nfx4L9z
Y1n4F+IZs5hSlM+RwhT7v8i7iFcHodRyQNJ+N1ju1C6qQlfQtsy4G1RqfX/sgYupM8BUI7YxIr+8
Z8RMpLvYDq2WJ7gkc7mIv0M58Fd20oHqG1djZ5zr6FAj70a4WvsI8C6i24eagdsb9V8L1XxHYb/d
X2BzKsRNdwIWsDKVZDNtJvE2LRCsmI1yLzj4sBsLYMwwr/q0bwFpSGdJO9y+jRhbbn3iZsnX60BX
WATbQ9hv4/nzwtgMj1j9uSHj8SSqSK6T2SbxoU2h+wFEeEnZpGEMSXTAlnVQhgN7SACZmzi3XeKg
Qs2XajQ0fmlmpHU+CvOHvf6gwf98dAUIhXRyod8QGa4W3Cq/p0wjbAsBvqbSrnx/DKfi0i3lW22a
CGRtjxCr40TSvktuGI+xM9zv/1QSWXXvufrRm4qw2zvmDmwVfZUYs5oL83qxHDQ6iZeadK/e1/hR
Kx9B+1XOv4t8HZRNnr+6btwh1GLyjkcbY2QaO7grA8cGdOQHmU3iRCu28O2MH2h4fSSPBonRrLl8
u/jsobVkwpNFLC4HJe0D+cbtK+ufQqbijjFgEbfdi2LFAQDgg78osFT7PXFQHX6fHsn4HMfUzx4v
VeVECFW/Ey+L96Kt82OpX5LlsgdSNkxUitIWfF8rkVe6IRX1XIYg6+32bZxrDy2lqt7GdIGD0lUv
5BEbknUvr9oGxNTGjgB6KyAtUtKyD98uNjs8alOZc0po2ZXkmve/L3TBM+rSw6OX52sN82ZKNcqr
k66I34pKsGKB/W7Abq40BU+p0ijl4g4rDf+OSHlQMwKz+hivB6Rb1HVWlUaRkzOkG+f3DDYp98ua
8s6N6MHZcqM5Fg4iaxb2WC8krfE6PF3s1AHRvHUuNUdCZfq0+tRyNOTr5WydzbjZLLZy+5LkgmHl
S1W3ZZUg/8QhNRO2pcKD0H5V5abohbFDfljK5xnOkJICYH7gjQLVsQcb7Q6byK/1pbiZX3jMLcqd
faDw6ynDsDwzqaxKBqDCLO145BWFCCRm011+oU3/5eHmaMmfAEINJx551XoOt/mfm6hW2d12rBzJ
bKNAYNkp9ofyjPU/Lik5ixX62VVzQWIm+oszgcXdzFT17fwDVC2ljBtu6uWuNpBVJZ9+nCr/f5g7
IoH0OKIIPyPVHLZBFDhN8mkEJtVK7sDONPyi5KN8YfE9cYn6PJho0b/3qZj77TtQ4587ay9Gz50I
M+CwwAC4/fDBkiZMICwgomLUkqQMCoOY37moGsxf2M1HcUvjA3HaYOLGjdXSFaPU1ZQiXiy2NLUf
kIqNhcTS51YWKVTZzHlvTOD2TxMlzAKLBrMvaIeYb5f/vC6ZYUQhZ1EzbUYTEHjEtWQyJ+b7NLFi
2AfAxCFAuF13bQWMOH+TR4rO7lCggpjETqF5EoK314mig04TDMHcOLgMOenSqRhxfWsRvAAtLbEU
7dF7xLmMI8DypoHFzTq47uvYNZ574cXqajfsgvOtWP/+BV1UsHKfXoPzSG2nNSLvTaQ2YV5CXuxq
n7IxEZledupCip5+YUC9csKOtgyzUt1y1JlZykWFruObTo636/uYOlp8p7mQCOvcnahEDBKbURYK
FdEID4Q3f4OojwAz1Whv1qYFHenpV4f68uJLRKJ/F2E6eE1v42nfMbOpzizL7vDEbdNqjXIC7wqf
9zk0MNO09WRmBnM+UtLLnQ+JkkpkFOf2YbXCVyJPf5VMAT4xPmcc+2ZBGMuWI7bHAUgu2nZhU96q
s0uq3mnjDoQO5so90t+S848UIL1/q438cJFqGu2PPhw4TasaW3GG/IUvDj8Ri7BvYn0iDNPy7HTX
0hI6s0iT3l+QCRMcDzMUg1BS3ioAMeWZ3FWF/LamX+qZfNc9eRVe36Jxw6Y6x9Yc//5rKlXa9f1P
oq1AZplMrnIycbNFilm+QoiFuJPO3Hg3VdPC2HyQRvak/M7Th2H5sZRVrPFeZq7V5TyTOiFV9jCW
Pvy6VGhV84G4IZ0dvjKIkbKmB/CDbCBYqAh08Wxm0zwrGu6NYsWaJL8Y8paXKtXiEi0omHYxGqxH
X0Yh6AXybdNfV0kXFQMu8BqdTc9OWyEonZ1TeU3OW5LXggcHFh+GC8Jqs1ncbHNZZoq9aHesB5pw
Hi2fSBIbK38O6ZDmTVcu1+vCQ0vUznRsRP/EzbukD7NwLhQEiBidDb63vunkRdXKCWq2OiWJOuc7
3npwNJ8tjC4hyD/zlBuBIkGhPneo7pbzfNSPc7cixEXCHNAcnp4JpHTds2Ko5fM+pNCy+zLsvoFV
/MwS3QNW7wY3RfZmvvfGFjcmN54JFicTrDhb9S7051BTONoPYcEZ8MOz5pQO8UwvtOd6jpvS4Zmx
VSFw8GWRX5j6xXJ/Arj2/o72N+EgVHNkj0yDn9dmaTTEZ54DkbzyZTQnOdtL34qxF0RPmVaUNgZM
MnZziPjOUckjjZCSIPFl9xxhPvHlK0aCqQSGxJzsroV+0jxhJXUiGipUl1tpvSPs/l2TDLc9m95a
Ecxo1xvja8T8YcxfWtNctjSav53aHkOjnLQexUv5ZGz+NYvYDIOfJt9iptXizy5lAGflfGi2hlO5
GUkptm5/0fwAMPNhlItuHA2Nbjb8B9BJYfLs5bVLDZUTiGpBcYY6a7aMj7IPfsDzmKf6m7Umbqa0
Xz6tKldsOqhVSET+B5lraaoco+2m3iD2Vf+qDOFxM+yNe4TBdiuiTifPhI4+7d+ABaqL6Nc1t/Hs
J9IbbmT4o8h6c4bgiFnjhAMJyUDgWxV+8aIzzsAvfoSUSo8BsKDSml32diDi7oau3EetmPy3IpA0
Fh/TbH8KdicAaQDaz4UnSpbZnYcOLT+9zqemylGZv4YX2EHv1rbaeJjXJ1mcIePjhCzLumOcY92d
4b0v1TyGHfDZzBy2L4TPzU8wcj0seUYaac3HHJx3pv+hTnZae3askoHiMy9QAnHurb86a6ObNYIU
eLKs0wgi3jAVO1J1f2ctEz0I8QW0VA23zbbH+KAuaq899N6lpoGP2IJZK8jJcE564gm0fGOZEBwr
AfgVnVNa2wzYm3NncDi5U452CvvpHJcu0ug8AKiIDUp90W4woqiO7xm8AqsaP5D0Rm8R83oWVmON
Fx6UheE+HGk+GoAJvwZQXY+yrzpfKORFlEoGJoBnudT0tuzUpbABoXz+o7V3A9oa3GDkq58lVAhu
c+IsN3grdf6+MBVlnCqfNz6Pn7zKjibES//zOkgNWhsVV9YyN1kXjF0sEMT3ZA5RthD0a/G1hfnp
VyCKLni0GOCJgTg3K6l1U8/Kt8bSBvD1yGNF5QQ8STVkCyR/lIEwueZN8LVUx49YMebyctGbrfv4
wMn1p3RtoBTWv+tkOJKm6c3AoFSGrtS/3WftPbXAw45HRC5nl6G2fygYrrFJEznyNXd59SivVKA6
u/ppmP1haJWN3/GckbSzJOmXltmtl2kGX2yX0M9lRhskGdN39GC/TMoVaITXIIkNnIWXkwWEjjBi
6qy1h2Juv7KVHxNX8P32b622ct6c79TKSxyzd/OrNydOCfpN+dFxq+hnTylyqp6qhgOOuxL8SP5q
XMg1qfACeWFXtTzSfjNJPpNeeie2Rdlt8NwTJi+FCXx31N6NGemmhthWXBevxZYocEwjpCG4pIAQ
wMV25VvICcKoqFFDYy9yzTdYZG7Yobxhtp+xpG/6MwAvD3kxVYpBRyKfyFKdfmST1DOu3TgGrbwC
xni93MatLLtw49Bk/QvF4EPcmIGjkZeIz+2dsNbZoDOshgUosL9G+l9cDxYSq2FawQtvR3fXhuVY
idazyBuQy9aUdZKFuUm4lJO6zjs3eyza3VRgnxzOO9TkHw5bu+ykvb834NhgJlRKre2kkLB51qaM
MaRRODlPuy/4DUyGVvMu4g1KMtJec4eEZOGqXoejfVAcc4NoqXazAOXRqbBLFS2U0ppLq/QTBGeS
c2g/R2iRpoldWf5k/N1Q5PGTVxQA77XwlP3pdK6KHeMKhxWBYCiX7YL+MHP7MRK3jQldZKJnT+Tl
S0TQGsKynKiCjQs4TV3SYKCgC56A0cJmBeNUt45cEmGTO17be0ejVfkE98/OFxw80xUvQCBrNYqu
zPwNHrwDZYZ+BzuNOxnd1b64VB6thfk5Atrd/Het4Bkt+7Gpqfenn1GyEzJ9XUnna+DYX/OfGqyM
9JNQpkSmtoRJlBmX4y0u39h2xw3b7Z1Lq1EC+nk7VHZ4CMox56nUZaUoKgD7s7FeD3j5u/v8KS7a
2PY+BpV+5c1kdsMadLXviltu2QIyQeD3q9NDiTSADy84Cmchh0KpzA4uViQEAnoDCdAL1+IIjLI7
HEx0gDvAuM8bo4Xb+LPBHADfavE5V+wwus3PXvg5rdpunBfrZtI7sIFbaoARABQ7UgwTwAiDfnch
ZuVcKHNtyC7j7umEj1ahfjvTiwnT40fw5rvn538mlRTx3LgG5paSRkDqB2YDh2bMntbMu+lFeUiR
7kJ1o4n17XixmB7INC7ZBVkokrQ55uLhVOkKcTCuqQQGZkIsAPc0TryrbPINXb9dvt7Jrtaw9gXz
QMA8sB8DKgzz+7Tkz2LuXxhSnEmVa59BWyYTj+w2sTeKq7Vl4a0XQFB0Y210YYzQyxv+F1c+9v7L
Ajg0JmAunOdQt32s3AJUgzcjVfIjez54toYqK8iZLcqB/qM6nIi4Wiw8W8ZqBLC1vV5SstCk5eyH
GX66qyA6aPtOgHRWGtYqAT0Nj/qwb1PNic00XaNtTXHTuZw6Darz9XqwHL8Mbq1m5Wk90mSPvn1b
7u5s37RehyXzxt6Ky8UBnlGylMb1CxRatGYByHDae/pOleApCr1Uh/a2us7NcTzfPmIbsQDSTVvD
dFehoA6iwwMotOIYrfDaYsxxXVGVzCpfx3i3m2czWeZ7i4ifeMv/fAiJImLggHVeoK+4u0uBmecG
RGujYj2lRHN9dSmDn9+nnBz09lV5syYWUL0yC/ENVuimpalnEN8GSN6aGLHXjPCiUx6LTZHFS9z9
N5blUUiyXY9JUoxjqCiXWDfvX6O1u8bcO3nZrE0f2WNsOAh53aZXo7cI3XeT5u2+ua5QYRKJ5UP3
eoBdMJJYU+KIxW3UrQfmSlPTizJNaD6t0VYsKg2jK1ZxR9gtX7ISbmFHryDNpRh9izyfXQS++eJl
0/Wbsr0UnOH0L+bXqe90o1JzQJVmqScFRU8TomC/BaarptuBoFY3tM3WXnFFsaoFniRU086Q+0lC
SEPdNF42OD3TpZRBXMKGpLRPBtKR9kEu1ICGOlIBkca+J/n9VhsXPWdr+T8YknJcZTZeEa/Ahqv7
KJXxgAiMwZjkWyVSLyXourwpINrSvPZksL3hWUIFtZwejqrYM2dz+n+ZG6Bp6BDvOBlxyLyfJK/7
eAQyj2DVJzuLL26UIFMTtkC6t8vE3GStXvMR1GrpfGpWIAqixegpd3g16NEZ47AlVx/6BS3sX76X
h92qX+eU+jugCKUF1DR8HU28nQHdQsrfbG5aYQXbj6R5ytJbklW5vBxvEeFL5Am1/RzjfOpMe2Pa
+pQCwRexSSZnq5rfIRcweYaVcR8Qu4xkFVAHbkMi4uScrOD0IyDpdEGRwuVXpsVQG9ycz3jBzT5t
oF36yfdEW1cD7dKk2K+wNqa9ouDh/JX0uarz6yqQr3PHNO65SvMacciwQVVSQctoJhLZZk5W3WhK
pQusAMLp9J86z4DYlKZaMaRWQL4uzUf6SIcHlGvzTr+CIySifpobx2YoR+0t6/cgXaEYCCHEmInt
UBdDVoauVeFX2CtdPLecmKAJenqlHaC+2mIssr6Bp5pzMT0Kuz1yzUQywswqJym+nm6AiIwFR7c1
lwUbIQyho42NOqCJxcGHz2mbv/+TwlEnDthnqIufH/EM8v0AlqfItqYludT0Qt9yhoR3RyKljQ+L
8srOQX8scFTFduvB4jTndLl9HXlzc27L5KNVuAZhLHlVQXyGerGYZeNqQuhrCQP1HVnQpaqm9TzI
iUc6N1c2RFMbEKgyHQ4qeN6g+7qr9R6SoPymefaXMi4wVP+/bJrhVeojjAud9EulP+Hwfw1rrcmu
W79d3hIjo1VjZRahrr45orXVzyq+9Kq9UlxhUPQbE6wqqt19SSXFCpUDQJEl6mnRbgzojaYEC1tT
PJqHGJURQRWr9VGEAazSIoJpGKwDRufJYrddQSCFYmRBmaWM9iKLHuVe9vZ1mzyAy70dfZgHjgpX
NmnFqIrXCmKXzwhLxvJwXMIxfWZ+zoebIFtSx01x6UsSJCEr22Mvmhn9XAsawXCFVWSF8/ZBTkBa
6/jQpJeA1E5mbEcRbs7w4CljiFqXXEuCUlMAalltmyxPFwPrLiZk9B1+ZOpqF80LMtX9QtU6/g7I
ckoJJCw4WxUhczyjXuKU1F4UL08cDVAVW4us0IdOTA6ovZmrJI+LbegSxIj5lTiRS4IEO8gUw1jS
m0ZHAuV6VkE3GDdVkq/Pa102V/eRkSgjb24vYk1k0H7cv+0mQkTiY21KIqO5mPQgMR6SuGyWOnOu
q0/7/ul44IBBTrRhXmPhdFjt0gI26VZ2dowXzxbntkjBB5ksSCaFBdflpZNa4aXnOv9jhzVFdV4b
sypdZILa9xbzI9e1+V6f3FUZkUsaXIAIhl+3O3g+cvjcTs2wXLBZKM3zUK59XE/7UFnN4xp7TIkf
IT473SuVvhDQ4pZjBHPBLU7gxzKQJeFC95aVSg7cHL71wO/02avJwu1v5VKKrfBEaLtQLLHzDO4m
5OaIWweekseRdWyspo05QXETo/GbjqxpILLEBx1gI2ff6dX288fnqe3++Iy2GGlqFhDo9YC+99XP
lPqMW1KpQ5O5VpngtYFdeooS3S5GOdTjr67+He0m8rJy6c0CajdXw6MCv9mzWG09q37Ax8iwrMg2
q0xVgJQUrGOLqwsSTe0O7vwmCMKdKETc+3Nz9Nx+ih+qLIF661eNJgvcdGS6wmMiM1n5cWFG3IX9
uq3s00uLfQd6bHH5v9Nnrm8wH47YRBQgtOgJ06kDVS1e4y+NgVUTmClKPBlHvic79qD/GHAY7zLO
Cmj1mf8K9OArxaO4WSNkL3MfoyZEbqr6vFKQSeCVxR/tPgIMvAQgM8aNBLYWlkIuznsPLHiKQqbJ
Diw7VG1HlW8kumtdcNcSUvao/uqQYyanWxW7wxxC881O92ax3vyRoUM9g/8pobYtzaAqHnjxq1wR
Z943OMqhaYjFktuG1xueISYmVLNNO6spm3bhQqTe0UQEmic1F1ezyXzJXtnhmy66aGMd+5HLYFgg
tWbqAmRoOFAxGKLwMzuNLGijTYeFNQSGU+rBYxKUZUgFA7VH0qAQEN8OMu1SNQP+dYxCZjIGQl8B
F9YO/9Nb+87LkpYY0sRKTvNGxODPXdRBXiGD+7KsxF9+IfjjkIGIwy13zhp4weE/qNHdAYJqVP/d
79e3vEU+p+ZtCDVvet6VnGGh0U1Rig2GvEqFHzX6RkHSjh335AgCXXFvDPYRMjNeakPRG/6Z4g9g
jO8rKi3RT5aLqs3IR3+lEM8Au7v1zIjXdBeBxbPX9s5NVtCaSaonk9GiPmokHsWqHWOvu8lAwiqx
9X6HVfyZHB1faM4zNenjGW4MVU6EN7ns3yeHIm+/22wXy8PStwhOtXvvY9Z+5I8PYK5HuY5WYq66
Ov54Zx55FIrfHswk0/laSzygIy0+E0Itqy55+NMwEESSwEyigFC7ysY1ZGtB2IvjMCNcCC+jp5aq
xL7FaOFhy3FtD/2Pbvd5LlAACSP/VeTAa7xf+vXyRI4e/e0gchd+BMVnM5iIalwANQ8QT7TMRu8G
fiH6b1pahnvgKOO3ECI5ZWd7t5bb3QCTy8XI8AOp1Dv9aBEdHXDjfMt5ql1Eh5vf9UU1iDg+bCra
pY+NeDyK6JgNn52dTu2hLFIFKQJxQtFoXlF82cAgpIdqiEQB4oAx7uuhxzHI1V24zpZ9WxmZKdH+
gJfYebNijCEFocpIDB8y6+zzxPyfi4+a+scJaI/t28XSo1IbBBJ+ZK3BlQYHn4y5m4rjFVg6tMSm
4nuRNGZ21C4wtRyQ9Wp3QS+Soy3eak6Og9qi1A/cMP7oAygoZGJ5uu+C74WuC+/j02CILZCoxGPl
+tx2biOiC/v57gNBO3V28uC+9xYkxNtcHyeJYkhkLl8MojWRdYNgJ50tAYQTOIBaMII+kLhr3nUw
jjlfHPEgw/dIG1KcsSIyfF0hCnKr3LAD5UbnGAXvKpIkSMqLFBI02C5y7Ns2lHwkmZZ+Dfpm3URU
yDDFiWWax4412G8LUAAHCpE8XT0/MmlVQi0NBLWgA4DjP0f8k5cOX8wmJpBD4yNRhEjNXZjhYVCv
poT9sj9EK+hbUqtJc8CE2ZUB4ScY/CNMYNL3+tU+mHzNqfGtzibg6O3YaPsjRiRg0Y7C4zBB5zzZ
s9p5liVycj7PIw2pYz0cmuheezfIEF0J8w/Heh4usLg09EwMr2+L+WoGjRRT9jeckgZJUbWEe9X0
EnMGDxx+JAUqbk1ObIoEMBHxxMNW1cq0uCwPJj64u7tuDkoYEpd59l1nMbpHYVVVcuA8Mm5MgAK8
Eg7Q3jTu/BEq8Dpr0bViH5uzdi3mqA9rRVUUtw+Psoh72j8K3Rgv6mVnvfaQddmI1AS8gHqB2Yvs
at5CGsBvgBnMmuqPW8t817obGfy8nWD8Q93mTG7U3LaGkyuMRnhhy/2/hZo8eUbgi6O6OGfo1BWE
QpXdU1QMwNB+ViHr78GbMMkoZfBk/JBN3O3e59xsoBDOaWDG/ZPWmpKA257MPcaMCG0DOhwfCbGG
fRNMpRRu6lb19xKEijg65nwzzhz24eJRpDj6xvSxJQGtjBmGbI078UYHkdh3bBCdyoLFbV6il2gu
ty0F4ZYsi/hsE2n4u/KgK7xfm1zbYUOkEUsTupWbvooZPAgIiCtBy2fId0QKCAqn4tBZFh+pJ2Ba
1ES+uS6tTSKmoXaI8bSPY6qZL726qbc06ZO0/+enTFhMlpreyULOKaH212cITA8TNbctqJctHvyB
UTDrD5D1aCKcZrxNAlOFeVF63gyVrffZZDTqUsrLvCDMwZ7pXyPyRmwQpCxIWz5nWuV/Ob4sZHPb
ZWZU9bYL2UlerRVHGRybR2BqJpPA2awEW6R+EGOagi5CKAKc0+DZdrNIZ4HWYlfYXqXhudUKMTYl
dXXxkjjZXLDM2tmlHAvf8w/KiL/9OCdTlGNCSag0QVXJH2U+FLzEIsfm0+8KahmX047qWIJxPN0G
ORuoAOkRkgMdjafoyfwJKjclV5egXD2znL1LU0akKXmRU8aq5Ow/SBGiI3Pl62Es2gIBDffBdAeu
eeffUtkwx+osQUzjC9jD0fss/hbxn06kozXk3DXFuhWFmoFIvL1B78oMX5bcXL18aiofX7OONhzn
XWAGWX6dbLIutOviLkXtYZJYIDsWJmmKkJ7mIR/+ZQe87mdTFHg5D8wbnIDHi3Zv1+GFmne3dN0J
xpLiD6KKSwgYeboXHejVSvIZgOhfnho6AmBj2bCHYb4W5HJPUDrz/hCWyxezlpf0P9uz4JvI6urH
2XJp5Q61LUPDvzb+3RKU5MmHDQGuTTOZDP8RHTxg+EKdtoZEDskrpMFIHPzlXYwtteRjNdegGXzJ
cYu5ufz5U67nMXr+ozXpi5Qy10SPg+50GJkbxxUKz4yqsVHICvb+RkNtKWgKu/DrrJIf7FMt3Ral
h+XPrLRm869xlkElS9xacBNAwFDPDkt+k03v/Elx2NdnI0iBYbP1h2KVzzK7XxNodn/4F1mTLbOo
PyESajqRt0EQKie/p+/Tebxx2ZRYE9lzXuaU9BaZHiHsMInHCrTZrk5/yZeCnc8Nl9KUo/9kGkwd
rOueluuwFxZ+S2z1oP+6w4/d3VYXl26ik9L3kpBk4Bl+wmssnBbD0rt3qH3wCyJl9rHauCSGrT39
w7Vado+RXTXYwNjoBgeM8JeyxNJ2R/wbYz8rn9UfPLVWFYIxMuH4fnPwlQmfBoo3z2w6aKj679TR
sfn1pmhnMQvAwEBp2W9BPe1DNlsgHPEOOF/J2wITXHEqRCZeDy1Hf1fEX3GcvLf1iskqzb/K6qfA
Fs132RAZ/uXrX7Bvg+5jRmN7QSY40heUqltH1A/UIfTKSgjeTnBdFFUj1e6CSma948V6zTrzKVd0
KB6pJhiiy2RQEWyNzxVT1Ay9WSJGGiVRcP3Z3nxLxwRiLC+rPuJdn4n9AGYCBMY04AwY36rrewDQ
1LEh64QddD3UeDdmMwCH0N8ljO6nafaPtmQoZAwFOkebcv2vdRXOLFmTU757xTXihjmgaDem0Bag
w/PZGnIE+Fc0ZFk4BsrGgkCcLiXsto5WiA6ZJQUf5Vq7ZsN1spo7kVThRApsHLxzf1LcR2t+v3WA
c4wG6OPJgy+eoXG3ouuQbpRw7nYmPEKAV8G1bucf4LyvMKeNvVIpuHj02A2EXzLtq+Q9TbdV2URx
tbAzkg8Kizh0aC5fXvN+tTwGmJm3sl81W6Q6gueOomRmVSWVHm09H+brqd2dFQCybBD0DTThYK0g
YLcU+tkKmZkrwLU582smqqP+MKCQGKyTk91TMnd5zxSKNmjRCN7WQPVdKjkzjJ7Z+8MyQfG1pZcY
koTF6xD3v4R0lCSvbS8LDEADscKEqa93WEJTF+l+RAjNP0TNhfhvRNmdoYGtPBfhyf+mX3vmLB+y
ptiZg5B78fGBto9o0Ox+kHgKqhMPZFuKMlQHgPPYG2ahdV4m+QBbnVWnrde+3Ad3YF48OwKzlBmy
hcf4451gEBHjnDpBcjrW9rzxzafmjlsg9Ztx287mSCWVTLsM49ACpvs4Vwe0gs8Dwrph4+zKIv6S
DnWfJkq7erGeSkokuJppX7y36lN5Tv0ScRDoQy5Qdt5uQe2xCmbwMMxIx6nWjeHUbN4skXv1xuZx
VIzKI6w6p6Jicni5VDaL4fqKkl0SveHxu934+ibQy2pTvvwBQsocdNXnyM7STNEIji1fGRs0h5RA
zNBZ+GUzuXPARE4wXdE90hb/RMzV/kUN/Y/NslQ4K10h+smHZ96/2ev/xiHBoWyhP/2cN4RfeoyT
bY+ueHiAdbJDJ0Kub6+9kKWquKho3OOqYr8UmxFw3QBBG8veSzAXWz03PXJ7mKTpz8q+0QpNv5/R
zxkwZv9HdXtKFRtRriykF0EErWK5Ne08HrOyVSl6OrXS3oDEcoZqBNoLYDMhGRmQCTKCbsj+wtDb
x1Dk5Im1u6wVSp3Zs6tS9Oz61lUCaQIkaLHgm/4cSzQlOgVI9FLZV4DmOWv/4AtVI4wohpODW+7f
O74fAaal8DpvwKyLQ5gWOIcbx8VG3xHY2QSpfDurHs91WlR4qLC6API46cnYKBBLxQfVuwD5GZ+X
u2pkfcqSr/2kjFdXCVPtrDu3Uz6iQU/FsuZulXBiFWHdYBJ59KllRYyKiK4ZcmUbh0C0EKpF6SVn
0fRjbexwXpywLbdrAt2z/lLIJNi1CsSAR1Lg61MYBtbthOdmbdT4BOiZKqcp+tGf+xBzdlxGgCF0
0nbgmU9JBqiZzIXCxy2BBqsdLBKeO6p3CmB6wXxQBRWypg/GSPEKdWSuE3dp+PXgNHYYoM8XummK
pYnxb3XlBxsrsI1cyfonPX+h2IJZzFAD6Pzuy8gDl4ZSE4p2vBWIuGfj04Tfsv0OEGuSLuP4ttld
wzzJ804elSanbIgwmtr1Cq83SUmd36PNP/9oZmZG4xxf9LQMRunqu4PPujLFwW+FMhShcXXJVZGA
VXlAme3jAUPco3SZBhyoCeSgykYiDniWZEGoOkdSpeXDu0ao0RbcfBLF3AoAI3RP1iYixt9fvYaQ
lnxwRHHex7hDleBvy27eVVbxqMa+QTGPREBLRXTqZJ79BlePBsfIricja8I7Z3YpINRjbyyEpYMA
affJZ8d+6iegrymRXCLaN9w0soqm7ZDZ5z3yID47cBFf2iaYAKhEUKQdIyDAclL9bOIDIPQbPjNT
t7WDW9AsEjpAWAsqRbDaLf3kC26FQyArUun+hoXwMFjMSWQegwO4qxh+wBlcwCfWnP3XqPtworb2
omqMV+1V0SrGX+wM0gYOugIe7yGDUQM48+5oSwDT+jbxXChW8LVUVrdTrnP7di0oHz87/G5QjNWG
Tq9XUgyA5tMhJBpUvb2wqWNXBVaEyiGfFJJP8VIr3z8G5Lp68szMB/UtbUPebkLavUTjXb0ymZbC
cgoWXEMB4l7ICJ7HckBbytwRXUZMsKue0zXa+KfcYdknCr7fIAs7vg+wTZAnkawnnmtMhUdiwEC7
hztMHb/O8GCEKvrT7odLXOb19PAHZjxCnx5yRVrnvfI4wvWV06NM79fAlnw31JkBN3DdGkmo4wJj
T1Z/Z+8ogL7uCQijm2b4IbiC494D4G+lAcDtPMQQMBl+2wyjKvw9HTadkpihpsjeQys7v0kNDGHa
2e8e3EbAj4dLpk1+/5SR3z3G8BbBdWGnYwFOGoa567VSEBZ6XIrrLD8frIVKntajPeIuifzYUkLt
XkZFt2s0QwTMxgw3ZAaVIWbJh3SFWTVzUByxorY/FfCiwPVHzr9Z7rv7wR5EpydI0jMDbiUi6imC
144GH+ZZiY7WP6eOrOApXefsaPjuRYn1TnLRf3xqfBycDXbdo7SBZC0fxJqFKe8N096ltUnwpZ2E
e3u8cPfFaEs2w2fxiBwezhMXoEQdPR4Rzyc1hr8o8/8djln4w9FeH3PY+AnH9zsPC4ZgQrL1zp/r
ULdH+RHBpgzmMmKcj9rYhgIMNtGVzeu3PrddXhmPLt91qu7BCxcbUExiK/MFqiNT3WWseBPdjtAP
waHTDEd1L124Kn/xEDn/JElA7spov9fpOYfCQrdDGiP5YPychyAnQvheI0mhB8wQY3Jj9x4OJrS3
1vaZ2RtKExuJNvBJxaFXApHqPp86dsuIuIJIkPO+lExJ6nL6L+hLYK7fpSbenMPRI3TddCU1RssU
ZBjI+2fWUFU8qH0Skm5+y5eG1VSHWNF5ipMkLUKhuqTRCtxIOr3oUXD9LEzFqkvqidXu5ydyNaYt
TcCPTkcxySKmrUoTSz8tB/joQcDXzPIB8RZqBm7rXzfAFSdkzPT0ghyQBAjYWXXH9KR6Wiuv7n2W
nCuaOJGxo2OeISNh+lbsbTu0cnMvzPSLrYGgNKg5s5ujmEGx/y/u97jRle6PMXfbzx+21/gwNrSl
ecoUPvpLdcbT4hv6BhiqAHlRuWGGa2ggCH95tnxCxn33h/U+1AQI/gBIhgHERvNipL1Bqb/PI2cK
aGvdHBLlHUcHW3dS7QxQOUW4wZ5Xg0P9BhEB2yC208gxVSLl/hKBYxGC+kQn3lQotKzZUIKBeh+O
kab/XNiH2s/hdIP/pSDIBbkv5hRb5th20fJbSxx9VbN0xrLlE08qyntcx6YJHqwI4uv5EwoumHTQ
obVc9Ky4wpJ+rvehwLQ+wkRVY5pEIczavueodaiFb1DZAcOlPYu/fizyrOOxJcWf4cMD5+p3MmQo
LD2br2QQwHpFOUb4iPOwsgSYpJQTn3nSywRHt3txmI0p6IzPmkuRAd5sTJoAQbs+ZgNpu1DaEF1W
wzw3vkwj6US0v9X+jHR8k9QvrxKsuZJIABbIsGi+W5v+ptpdU2qsMZj/UwLh8L7zrDUs85eUx8r5
EsPR6AchgrqZuXZgEWdObsonEmtctZIPjE2RXovYC2VNG/s4WkNYWoVQ8VZ6xXYzJqZXwBq8phIR
tZiH98WDrKI8I+w5y0+szW3DqKZoPVABlZm7p9Ilp4DBum2Ha4axYylM/Do6VJSXxg6B8gMiSvUc
Ngd3vYhIXgoR/QJKM9rPgGq6cymAtD88i2tc9cvcziHa11OxaD8zESv2VuJ2+tQQ1WCYVF8a4pcJ
FWkuoz7zE5g9G0b62F7SbC8zuqGXgHvPyXrxXEUhuhXnkNpvUh5YCzXBcu5gNXNLt2Q9WXvtq6IR
0Wt/Rn+4yvuC32Im4dQNBlHk8yXLlh4Gzj6fxYcR9pl2/ZUs+TlqoxL2GxdeQAgt+hJB02inmvWi
zDJtf1RjDvq230vs716xZ4QzlidZXil6JdlAuE8BtCIVO8BzkNmN8584dPWwSI7MNKWJ9wo191rD
1wTZdP+TZi82JsGSwhat9VO6v27jn2Ue3SUtzRebUQwNerdxjhC8N866C5XslrtHDp4n5Zv3AFtw
7zhYrN+EuUZ4PfoWpTlcyr1VMTd7Mech+TZtJs9hPKHIDRtzs0jKvNc1+oaOScbaOH1BMTEVr3/I
Mwqyzd9DeAzu+9VX/bIfafKRSX06d6+kVBapqOa2SAzObZ3jF+DjA74FPN3KeVnSzvb0nq6+WH16
BB+YAO3qi00Q8ULZML0VUYKZu+YybltUf/yh4TAt6vY2uy1ajPpdWt8n68dvO63ADZ6Qugg7W0/0
Ni4jdLKCvDK/iN6/lZFssgeW8VzhC18Vf2HoobzX15ILCJ03KmlWnyerj+/tC3CEJNloKyHR0NcH
tY9mIUGzC4OBVf2JClfycTUwo7A28BkOq+yGAwc07zce7bnbZipND9UxTcLSlba1+r09ezpJkrU4
InJ8nU2p4+LN5Oe32fdOuSoHi3QogTkUmwNsTuft9MMyiRpzfeEZ6kyboF3kcnKdVcDXObke9wr7
mdsDblbQNfCaBhDqoT2JjlbbZd7tLAoMU5yPM5T8bu1jqteEJxnnNY4zonyqjIUanv5+gMhdL0wa
jT0Zo++LaglNpmGcoj59BJrPtm2LZN2IIxdDAJPruY2gCT7i21yILQ8IpPoZ5EGDhdf2kfx/Z2cz
Fc6ZrJlUUbZnRs+1p26nsSmXEPuQcJtoilEDtqt2ETYZYicVYetJB8KOGF7m8GOoxy3FDojoK/eR
SI10FUIRg5iRv6Pvxyxh4EJ3G8vIzmXkGHWHwIvtpXv+tQVX9medLsPE10QLs9bSrqFgliafIBT4
ZdcGTe8MBRFVBKUG7+s3qIU9IywahCt+EVqWVGvsEnr0A64HlKnEsuca91sytfGexo+X+oPwrTRm
D9TaOnZUVzqdL56a5UwnY/aTuKYh4V+bC4OykYPg/WHHkGjI9ePikIt0cxm+Cctu9mX8M/ZrMlIm
X9jPQ45BaSG5zYeME15DsZ9PxOUXVaqKADtJc+1c/aFzE9ljYg6uJ7k3u2tbcykTRgt54Ii7Lb+T
GxqxNv2fRMP+87Y2YMHIVBe9fXFH9P1ixyYukOS0BFMiX2Ep90tjsXDX2QUCJEoakBF6twtFXWYS
+QfEJg+N/tCDRbrHrs/OAl+be1Ep+2/b5iNkO1ytyPQVIIEbML/upmx8q/mSaK73P17EuUQgvyD7
5DjefduA4KQiv9njF7n7MymQF07zDSyZR1pYGFCmYAtJYccKGZDAtS3C2olGhQNFoXLHlDVFqMJP
WC4F6l6Ajbnpa3scCVRmRANucwyiKo/oZvNOk09Cw3yQ01GjaPSdESIvCVqemSDGFQrubkmgyGEy
IMkjd+MEGuW7t9hiEgI3KNRMD8BRTqceiSkDAsX5MuI5JGGPUCJFWOj7dH9CUyStXw1RQR5bLGQG
VqBrQ7zQIw/IztdNp+S+1YFj/MlPw7SVhrEprb2CzaI3E42fU6iiFQZRKRGAhj9zdRkB8GD/RCbT
9nGUWgZCl8xqxVAyZcqMh18+nKbD+XRa+ysl8/muUeX1qWY7o1jH6Hf2+VlyCF3FIpUnqyI/N1ib
aCmWTy8yK/v2QjFxD+/yhxDNdM0a1sB6Tk77FYAlcHyXyh7UVFOPap1ZY4+cu3fq25ixOyr3mtmX
6wGbxXRh9Lvi0adNgRHX9uHORxGjzRxFCys+2BjoPiEMymcuaTacGXomrBkPYjTBqu5nlyoINIEz
/oHHFzzUUvJdmrlm841hVv0LYW0OVigVAfea4vE+T9+tZpA/4daSdCWNT4DisGZgbiJNM6unPAOQ
bSZaxQ2bxvdd05p8PjcQtjtC76px2ga4bv537KJGRJ3OCe1tWPyrDTvzLy4ALCGh3XyhPpkDhtGv
fjg5F9g/T8hTZLiS2VpQP/7UV/hs9GbJmX8lpIKF+5MdXRdCuJOK6FXvPH60szQheuAORizco3xe
RVcoHzUh8u19HDR4FNNUZcmZqeeUJic1slUh1E54pFfmJoGQ5eqbkdexUYwyM5+53p7WO2uvLXC4
0nvXX5k6ywC8fdxfEPij5LihHJknLJBSU+2xpqTahJ+QUtzS1k8J83AgMQ+B3mg9F4+OzHkiJFcr
jvIqXRJGjOlco6KqzYv1WZGH/iSa75Ig/XdWgFU/gSVTrf6/HssTjWYTucnD/sNyHRqDFj60Li+W
Y9KU6KQv2sO39KavVKNzrkmEUWr1n5CBhLAUQD+VfEm01Idv3PZpdhqV9fXDMubGpYvKNftbP61N
5uH7qFlevKcLAv4H8nmbTcb3OVu9QKfAxeUrXmmhhZ10WkQ+MLO3z3FpOKlhiOKTfhgeVduKgJdP
CcW00sli3oAejrO2Dht3dRXLtn3q5jpxuLWotNWoOvYiI4gJveLBQtl+//bmmfSSxqfO5Z2HNYdi
tQuFHCMnBoh4p1YsTcGdMMk7VpxuSR3Xqt+MBSU0V6diFmZTt7WMapkm1xmonYIQwBMKP5mOHvjJ
tgSdydj1Za/BY79zboBGJsV4UwfZ2suLN+ax5SPB6k6iNJm+Zz0TGu/kdrGf7gSm5Avi5Fj8Z4jd
qjZMM4eSCbTFMDBH++m+r03h90WLCVtiSkziVwjLHweMDIzJgArqiL3X6VTXa2pw1hA5bxO0mIx3
eMsFzaW2ua6kq2N+ryS7drmLq+/bdPp48XaokHI9k9yvDG/P2inX8JhrSNDRDKCoI9C18sMDyoOG
AAOG3Bhb+0zgmtvtzOahw9XHdOvFQkEEu2MraPDZIh7S8ZJ8+Q8UH+jw3e4LTRO9z2ro9VkPKVOd
TgKuPeAP2vBNesem2VqQbgKlKxw90T+qT2+UKAYBozSkyISE89IAyU0hWpFHgR2/qwiVeHc94ebs
AqSQamvCOgqpGP8uozySU8+3H7HkOf9mhRiAyh5rvSmSRQGBOPoxjOPH6Fzc/UGpHyrb7RvEOPux
/+7Abys18MdqWwhqNL5j6IiuTbKZXnzeHvI0PojuEKKcRh30KBvaIDw+H2sZwq9csUICvNIxydQ3
hzp5DtAZ0CeXii7bZzvfE4zmHZlILC7zN16u2ciVd1oYZBU2XHNA8B0aGBGa4jv7lBo5uwPcTMAE
eg5GtxsvS8/b8PJrCR0x2FZbG1DVNTPkr7lh8M8LnLJpBqqvGiAH6PVBgyBn099CQF3i3RyYQfQT
tsUw0lJ0p23j5F7pKKVJh5GwTyYfBrD7JPJfK8EPxkYehPf/PQcB58V4uAEY9A8LGDZ6GIxzZlKO
QjxfrPe6Ub572LhsS+CQgoT9iBrbfZey+g3X5Dorowd3m84Z7taaaVZdXKqhiMtjdfP3woNGJb0M
6kuz/IMB0WCOTiHBqI1G+ITENbBqKjqJeOh5QvDVTsRujI5O6veBeibcf/X2BqnMW3JiHWsDkCsJ
919IDa9v58KhBQu93uTzAtzPmJ3ldcd2WPwE/rstF4oilM6Tz9UPYdy54/nZQGLwiKd4qNklwr1o
EKGTGWzMsGtzmKtE2iLOYh+4wxycJ1/oHYZt2DhQZ2dKkUaZ2Kkw10DWBcIJnBACRBoSMawcs+3O
hARzi4ybFJOrqe6A0U2gmoPFTg5bbmiMTHtHRvsLb64iyW4PnDE6zjSopMNG0Hk6AusEPtZdLZvX
Ijep3jk2pRBo1AwaJrkACxtNzPIitqmIBqUqcb69HYXJLoMK5lhO6wZ9sQotuwET9XvLca4FiTGn
Oe7N0Llaba4L8+xvUp+CQ5dCbu2nVot60wziWm1NqDsPiwTARJQcnCnsPZ+ZGkDG+QuGpgEpSb69
5b0qOs0EYLTKYKdQCtnYBeIjnef/4Hr7mAH9fG8AuIe28UzW8qS1M9clSUpCrx+K+wWZ0Q9FFf4T
zuLsuBUssGLBtZ/zVA5ZlH/50Rj2nd+MtA83jNqnBRILqa5LJGWt3Blgr3ps1FiSMdnHKhIR7/eE
fn6SNpK7ikcQDliLjf1UYf/0X40AKtmInH+he2YBl1RTz/tpQXmThav7OEiwgUxjkW77uzkPGfFT
svo3tuuVDfpIbK4xrAKs2P2UhYQTDz2VKaSk0UqfTTVv7Q2bLYBKAxy3rAX6Oy3bFfU6loyORCe9
Jc6Qx8lZ7y3629u19ForZQOGqnEYGjBHeeD7B3GQtIAml679cZXiWq92+EDCBbv7rUZBLnaTJ1Z6
FuEI5ovphnOZzZHwR9utRsL9PisAdt4EtPSXGxf00uAXmRBb6TKifA+tN+0KGqDs0101x7WPoXjT
+cEUBednuxfJa8eSqooDTTgywKddq0qiD4E5K81sWjricx4JBNBAehTWVcJISJkHfikLIAkKyAbu
wvrYiBWIvc9dyiQQPxQgHnWuTnSqX4ncu7rdhQPcZA5Xc3/t9IJa8modqCZ7Scp5A/hMptn6tJ9H
F+Bt+nM5aRtFDAaLvv/XRqzznyZekurkT8hBLyoAMtFzj+1QunsZIggviz/KPEgZKj4n5fsgEl9w
A8fd/U+hRIZ+lJXszU1parJTrCJRMG7UEgiEfbUhwtVR/eTxzzbsI/y/xQT+dUAtsoZKQNYa1nOs
aC3cBim2F8TX2PfgyTauMwH4wnNvRTFHEsnzXiX11dZp3YRxe9FimkWDeJGLUbIrshIVj2JLOvCH
sPPm25VLv2TaSpdIesreM7WnRmxxnMa6vPOPVCl0bwxOwO45zzn0dFDPZ3QDLM8ykCT7ueCRnPsv
++guGLW1/6QB4fS5ud6OMagpCnOz2Z0wLQxqoYKXYVWeDwsSeEqKqFP8eYbQqEWlt4lFcBZ8zZga
e3VRPRZHIwCvwr3zqjuSxiR0k+2+mjwKhEehYTPgkjBHqBcHyDvqqZVWgzd5GQyQWsXlFSG5aLph
qgjy6U/t/nBjxT/65YyhGxejBwhcjYmWAn+bFtFQG4ktWw2KtXIo5vitpU+gFOnCJYZ4NjmmxA8G
Swtwgv3Lzj2oynKVmyY4+7C7iI2Y8/AqikTR0KojTwcRyLeBZLDZB+BmZNrKAUxh9ae15uSc8a1o
WDQvD5j6ocKhghicfoMMVQn5pfu4oCJKyIYMgwcgAZkRiiM1zPp8cJe+ykqxccNa0OttiyYt0CyN
v/HBpwWTsxzXTxfCYJaT3pS23emyUOzk6n7z+iQsJ+o0duR9zdImgtsGwmSyMEPwDeOWTZkn9J7P
VynInNwnt4BWJ2KUDDTsDLKHj4AWlgUKAoWJ8hkXH2KwgBLzfzhzd1M/iTmHw+twezmGz6Pgh1uw
63ngWvGQhEXGIprXFL1BDTafjE/iMu9UmLcXqspIpSn76tfmzZtlKVNEzoKIw49FZHVNIquYwaxe
d7s4HlNKvLOTNb2pb+9MMWyQJWH+5d04b+gdk0Lte2D4smjYXgPV6xoSNZ7phCeEwddriaALJ+jj
u5e/086iwf4L+v2yQpuk8w4B0RmBpRYB+yXsLQU8QQ5L7TjqbaBPDTYgOmJJx0BmhvDVu5ywRYcI
omiiHchP0Sgll9YzUHk9Ffv7vTI1/Nh3H0vsrAICQEW9jPBEnzA1IMLcsd+AusdWQanm4HZKwCEZ
cUzNgXM2inoqJq40V2B5HizoJOMUBLlQUOK9PKyPhev86R62O+uXry37jo8jC5QnpKOX0CiYDnf0
ag6o3FIzav57eYiJStARVhBTDjd8dXLak/89ervSn3lCU6JzsdvgMMq5JXGVTEV7WzTZb72aUeta
ljjbHlNUXPyKXYA2PqWD2SiGwoXHxBUjKx/8ImgdKzyx7pZ6+kmcyOENaYzX8QMre0x9bCYmPSW/
lTmfuPkQKBTOjwKrYS7PLXtWOdGIVlP2TYBTbmhQSKA1XDWqRYHBBRA6mYpHqq3mdhcudO8fHBJX
oUG3Wy49axoLkXIMLhVnuGbnteJsNYNbUxahRCsv0aurxs+1KoL09SkAblIpK+XxwXom43CqycyB
9wHwe/gkSfhLoRC/zUP2OBhfq78lQ1REkRVptGV82cyb1eTSd/3e+vPKNil1Y4srzQreWddod8vF
REXlhow3qQQQ0OCdwmxyUQXnCjwM57saLbmDPyw3M6Q4rrAp2NlWWDM39ZWm3017fdOPbyHcxEXO
tyT377To1VbI1HRadxlXq44NEhcyHney3mhG/nF97HroT8gHCLpsD09WL5k45C5rnzbfCPpsZO7Y
+QilIXqn555G2nRReiuhoEwPRwoAndL/dm8KZCwIqULdzQDq24RuhelzKxulJ5C2petlaAf1XAsP
0VRBhP0haU426JWu6zyo5yYauePuoEad2AW3HxXO+ETgtRWWX4jKrjcGFcM8VIKYjJpNPYtSOpYp
egWQRDfeWrxEY1QupT9eHGx4l5nBRnFFTsQQOIBVAcRc9tPf8ekbRoCVFeWbArG4JyrdoJGz2Tsc
zuBtSu+LIUjbsK37n8qhD8PO1I+w6Edd7CtyqqICQWzej/GKS7ux5J+WRXViswNQn+eEGA1fFk/D
j7hxsdWd8kDm/NOth/T49rXl8M4PvCy7i+OzsZOpsnbIaDk4ncAyuG24b82SjYdyl1k5cnz+QxdP
wkRQTDeN2mD/b9zo2ezG2RrfS6WSs2dz6t60tmOz3hXXBJkd7WC0DHy00fJj4rTVnFR3f04kSI+U
mN8IoVQ9NnL9tsPX4VOgVYmwbLHY/eia5OHZ4z/UM3wijpc1YMYaHskAyNSFtDMOBuuNZzy4jSDR
4xQxNe9X9tIZpzARyxlROQK31Lglx8yBEOWKM5H1WaX4B12P6UWnplPHYBFKJ7eA4jGjerbxCI3p
dJKJBXAixsfUuUflBYpzei3taLcig9BNphD3XyYroUTdbnj7Kgsbk0LvAT7UrzdVczosKux/bm2F
3TItDH0WmbxNE5ry6ne5bula/YXjHIhPWXwseNJ6YVYYlE9knC0luEjugnjESaVbe96VGLgydiT+
wUPlgTrEHRRmvu5R79tpDP5ZAZ6T7xg6XMDRPHlIF3+IKnGMrm102a873hLdsGXLjwk9I41ppHuI
Q+gP6kEEwe7AzyfZHz1yb/2G7HBRfGDW9nm/DMrVlMFRev6zSGFJIoBmzA6v/KMHpT7paea5J+oN
zHOQGS29juN77lK4kKBQO3CMzzmKa1vOPYG67JNG2W16BXgiYIFiHposn6nT60JKVojNO/8fefZV
7lEP5sSZdjEmkj1CeKdXFk2zn1zhP3/XyuzzJc1yCeKJb1F2QOvl/p9DDTkUxnTJG4a5DOUD/y6b
drbFgWND3+IwQvCpB3874vXhtFMfu5MkRIL7OS+rWX1DPXX+59aSd4UIME+b+RAY2Orx4wiIwWP5
58jX8SKc5zgx1wVqiaI6qCuN4mxTG98d6Q7vNF89UPJOYktqx1FOed67rxA7NpmcegoCguATCVMi
70H5PCQ86m6hIrvM7jJuYFUbyRx7gTO8qJ6AOvR8uFgDbpqUvbN77my5BVc9ke+rb8dTJgwrIRHv
OBqktHl2UiursEgzeWkSV6dFJ/0R1O/EbnjpX1EiMg56TSN9l5jOF+HggMB0146X+I80QEuidb6d
OH9N14I9HeLurGbN+KdB0rZTFtGB0FouB3jN+djPaZfmKA+HDpwWLdHvr4gPUoMUPqnqrbMdkC/+
JRh20m1Nl3PbOwXfpL7ckZITcRYBEQoL11APyD/+A/3TFoTgLdBXsKOXwoMU8IfPLtIeGk6b5m9+
hBNSAq1g7BJvqmA97tFmScaczNjShTau683wbWore+DolhbjU7xd6IQWrOCuxwkgwv7KFJG3XQNt
Ni3+6O8HkYC7FQaWGvVDW05kfnl0xMKY4kgoE8F9quxv0NJWVRZC4D1ii4pFSuTJvXOE/SbvCKxT
LhGLzYRvoUrQaiHhyaM0XqsmKR0/TKLig/c1nXfkwOjNwpXHIuL8V0sNkYTKJxE0WCcFaq8QPsWK
eDMeHoooBM0qxQrDZhGr620UjAexp3T7GH6XFZ5fY/MUJvOheXNMqKV1Nw9fWrF17WkngWPr3vt2
85/SiYGateIkyPFp9iONy7mpXJMsoRxN/JHQBMZGXe40inLUi2jAVRWPLDByA+JhB0MfaWTafpsC
ZNPYh8k/B4uRLwODw8AD3mXHfErURsosFDQFcqfiAtMrVT1oSt9q1gxK18R8PnvQtIdQv+59vTlr
B0R9YlGRThvWOyshkOeBO7I8wQkhi86gTYsjdLc2KD2n9yPzfTL0nVlJZFz7lGleTR18CQbH4Php
7bucHpyMYqjye4NJDFxePTqPdtAQmEGQ3HzpdTfnisipBUpIdxgQ9gEFdwOPy8lAydnQcsieRkyc
CwUd25+xlGgGSFkQ3ADSswpQevwtjR0v3QrlrpSFv9ORn2e+mwbqj4LmVSzv8n/UYL7VGznMhl9A
nFAYDVW0mmjZeWpy06WrHxXJxr7u4hC2HrATOxdZZRj04gotLQEvsTlgIrXdIvTXHU+NSEWwraPE
+TPl9afjbMWtkXyXpbcgxm8HQl1kxVMo69Gbw5ae7HBj241M2SIUlaMbIXCde87TwSFtB3dklg+5
pQnAgJp5Dt/bc4F64FDS6Fjl37c7UKq7/ahb28gzio2fxgZAxRGA/N2xT4n2E6DuE+OTXWavNb2C
mZBdHU2P5sWmgBr2osVuYWICSWXX3LjgpUMvEe/kN4R3m3sgWTj/8agt1k6nDokaef5IG+rmz7Jp
pP5Qn++dVReJWbGu7TKl0DwMfUD83BaUmPnXyxbYASv4to5iG9+5Smrb/dwuoPUr0XA/uJ+2MmQQ
z1Dts93crCKQew0uLftedIV8OfKNI/bdQKf8gW1HocAsYhpXQ1+r++O4MzxkewDdO5V3oQul745d
77uVLTxDXX5WSRn5Tf5LFCDbtHYZHm+TNFHLD1if4Rj/4eXAo9HMTlEBS++xC2j4Swg9e/yJBPvS
X52IgHAdfeZ48zOp+2iGw7uOXJMT5lFk+/FaMOiMGEy95VTpCYvh8RHDlC0JvoQArTL3CZTyvlPJ
edW0p5l89+O2oCV/fdtbSpPpJr0p5UjAnNm+8f3MOqT2rVTr2hwRAC4en3ZOYp6VgoS6pxZhlnHl
rGgBWezBCAokQfKcB0J/BOT+AzcFX3VlzHRTaWFfTf1fGV5nByWA9NsB7fixkMo9PeBD8ZiC6NvJ
ZjA8AMbRy+eg7op/U2C3MFMbuxxQ7yhrW6U5SQ3ssCv7zlNO601eOBUn/EsfHyHJZ5Qtp41+HwKo
sCvHScAJTvMx8Bh+iyF2QSRYTuvMGPMw9rJhbLZLSXtJQHdvAa0PmPOsw4bqDpHNvw0nahPypf5+
Yi/iIBvjmNA1mlp5DW+EvPyd8vmMaQmaTSYHPYYJmcItSgLjMGW2TxyESIEU9dQOjpQdjUrVlB5b
ZWAQtFSMMaC2Le9UpzOZN8/bCmtKUtQHWyGi6pcE7AISSrNMZ4zo8zJ5JvaUZ+oXAWw/lUtPPpYV
zbeWPXw6Yie73UD/BsazaSEXo6ltZsSMeD8xNrjd3Oa+ulVEN6YiE5TVFblT2gawoCXWsExz1xS8
ECKldNtwBJBgTsbLHNZrALii90CIHoSQ7HdJ0+uuwARgWJyu3f3leZfXyd8hGORnnqeaWuQJYYDM
1wRw0qDHC0GnFYmAFn4nQ8zSEJGBfPb2T84iopn1NSQjxxbZeojxTcSGYKz9BXom5cIlUd9KSoXt
gZA7SqiYDR5iZNfBPunUBp2Z46M9z+JffkhJ6/K2BKHiEbgCeZ/oPfsBQXYVtpUIdQb3JTKYze8z
DKDCHJiRczvY06a6sx/xV3ZdRw8QDu596xqq371q08/YYNh4jt+CGlxivKU3NdD86wlPzlT6iGV6
yvwqG5Dw0H2j9hnehfTHdbyqYasOShJgLLaUqdgQaLOhTuA/u5qeSa5EBDXib9nO9808B6cMWbO6
fLvbCevxNrKzK/IO8Wc+8WiAtQ1+uLiSdOsXE0JNSS7AQVNcyMvaiNkNQh+BXboOrMc2odnUPz7G
sNwBnZ/DLXTU0gNkVtxGqTIBfz6ZRCWaUFVicJOMpZ2xfMkkhf/2MyzRiqaz8nQmg4ySWyWw+evH
RqSZZmbjuvdlrv73zKjs+AgyGRY1jORexuQZ5fhJOj+GWJLSMPgVDJNwjhnhWHOIv3/WXe3BqiW3
BTzJ16uCpju4eHvSEFPCt09/W7KHs+XXO690wJzzbaZ6zcD/EISto5f0pZ5UrcXnPCHMpFCTbFoJ
/XAOQ22ltayLaHlhwtAl2RbVRbJOGoQo6FF5OwfPjM0jg9fzgO+WAFBwEVtBIaLZLTeMVKucKeZk
zoIYOX9vghHmeaYut2eD4RrcztDmYHYjNvsKivZryAVWTiJqwqJN2zbcqQv2DuRRmuPZGSQHJUOZ
WNBQmFAwmuioOVi4Kuc3iXH+ZVvtjIqJoGrTFwDflhqJzZNA6hCIpji6SQwYJHRNjvbkC0cZ44su
kYWu2oE121pkqGH+EpzYj1/4z9RnchJWIp5wzQ5ipT178T5i7YnwaZZItnSnIt5d+AraVnPXw/4A
KTbUrk62GOoFLt/NI4uVHrVKDU8W7WrRTL3KtbVCL3WuROtH8ooN+rdn5SmjNQeMWpvgjDdgXOwv
Sc88H1e6aSFcZv9Y8SEv5aGssdvMDqCxBFpuXxCEZzMwV5RwAmCcZMzsfW5zPynAfXQJ9M/4gB/W
Dqyq8psNXmGqwJSXWDYmNe9wNLsji6/V6uq3V0D0dULG9JjI3rHrd5dNy4otWbxQ1WmOX+9/1j2g
IwDRznV1BwoX5rcnk0zaFGeEIBPRKRNxznyJAAfXa45ghAgQCe7idEU0/Tv+Kg24JbP+XaWRfqMl
eedbBg+DZK8Hnqvyk/OJQgAFbgCqNdBOYRjiKR4OZHrYbkiwm/YpCeeTqP0Lm2jC7KJnzAOUjF/n
KH7+8nROhGnIGtDLCWRfGRJctPIAyMZtG4cG/AJMokDC7M+RaAy+A4Flte8brqB3Gs/nMxK1POle
9RjFUHWCaZ2up5DioVmHuaYrdqoZVF9+PSWmgMQgrL4lFFSnWONjAGMmqTGFQwKc4/2uhUWrGaNb
gUOivIb2biGTWpzb2bQ6sAWhsMJhjmu7MnB3I2RIO6Of4Bbh1EhHDV84psB/FrjIiLlHra1LSHdq
07WMGo0HuvvLMpB3SpHodzqM0fzeNKg1FWMbrAx5JIPNPmlb7CG35wTiKNJjR1nX+LPy/SOimuxQ
3Iz5GbAx1y8NEJOPCoyLoaQqnyI7J7RnYwFqNgE/fRUaKz3HMVAOciQgzYjP5S2PymnrRQUVvmtb
qjmNNWOk177468xayzp2+14aNnJKJ1zZJEYnHouRky2jjyxOGtyyI94s9mceXsTeThMNwluqFz9V
g8p7WdowZg7toKOY2yCVpwHc+giCn1BEHTFssQTkov6OKFn0jhTdqG/z6NoW8tHdEhD3VS4SOntv
uHnHeV+n0Kn3vo3GzF72WPgnOt+GXWfpPUqOV5O3Pe/eCdwuHxFaDtsRXCHONY5T9KwJT54q8MsZ
AEDb477XgcaYq9FqpB8/aEDR/c1EY7+M57v4zEs10lj3Gmap0OP1MzL3W5CGwXrWmQxds97VNTND
q1EgK2NAYgQ6lxRRwlPbuaFVv8pc1+HDCwKustRw7OHTED4iyZARm2m16cOh6T+6oQUtfhUI3B6o
mydDxtngwPXWWllEEboaDAtnRmEOM7BSM4AqvhaHoGo22st/e1FvRhhAHSJyi3eZFdFDYEw702w7
4JhjQA/32pxZyx7vit06eeMTs+PWc50SlEC4TxY5lPwN2AbhQiDwYRbfoyurXTJ4j0EvO0SAS1nL
aS9dvfDvBMEIdMlMfg7Fw5nbaJaY0MH5tQIl8tpi+6Tij/eowNfO7iQ3+JyCr3f6t7he6u9wVCe1
r6syOoi74mIKhwedORjzAOk2Es/p8I2kHEaG588XIdfffVp+f+4MaIeY1xDfWCfJ6qM0Km22afrK
PZJ7pskI2UiRFfe+SVAFa+OJCoj951kTuC6MbG6Qox3stuPNv/rAZSQ+32r7j+2hoBvf3lN529vp
7vC9SpSJYyp6qUW9/OibBudGekFvi5CWgAOJ1JsofjQlZNNOBXE1N2U+gc7/2U7gCrKmPWyoYGfH
v+sXqNYGYACsYNen4bFZzFEgFn2O9VXKjJj7Ch88/77IvqTj9en1vGuYOmOj6JvpewEaKZSeZcOa
5ziggSpEMd42eAkdNWFmxeN9Ut3vfdS/yW1yV6vzGNnV5X0t64JkvGcWWlo1KphJ79BnaSkRQLp8
Fy20+C2drGK4Rakx3moR2YguWJmi07nrq6yKWd44J7dDoO3sdIx2GTFl42gftlibVhz4rm4bTtB5
G8JfE/qRXqMtj3Uv5FAsbZS/hT3Ef83FbsiilZnn5M8HqFYYElpfOHB/mW/ar5hh9lvsQW5EhWn+
V7C8tWxaai6RkSMFm0iHDn0MdxzHi30Yrztroch0rVmv2WKSAmXy0o0b5ggdFHmuTyC+ZfP57I2O
kzBKjOsDJhQEEuDf0dp60bVN/AxHeVTLEY5J6Aw//q0CMQnY6M2bQrq67aHc5IDhN8O3Xq2iAgC0
mYUaLrvQeQjEdx3Dc938yN7l5SW4xSTksUHArWwW5VBD9jhbM8tQh9ZhTIsbzjmb8Kfh1K0shalJ
yCJugVGv0CO81lCry37j+a89AenK7uJ+qqflJeuaIMs3qiHzZtz+9ssLp4plAcOTgj52RebUXGKL
O6n3/pYGamFlAhHkCTWQ957c7rWGzwiAme97FFrsVRp7WB+0wvULuvGLOdRUb1jJ6DHMLIy3DHW/
hCabzuR8JdZeEIjN4xNQPr9BFdyqVSjvWDW+xDMQ4+qZun+fcYo0rFs9JQJFbdYuKYj1RrVVx2Vz
SprEZNlB7660vlmPGCo4pyt2T3ruhflTYu7SY0Da356Wff/+AaCrHmdRifxiOkbNS0VZT7EBJH6X
DDos05tad2MS873mrDKH8jlRHIHe/2PmvOIc4AtBSiX72GsdHfLef3QmcVUFkhfuHVPclkZ+qwgu
cAc0AkxUBwBeHQmTlYYOyzsW775HR0wZundj75hIyiypqcfhPAWgDLVvYk6Z2JuDUkGCypflrPsy
RU8+udnvVEGUhRbM3Ci64ZHN/L04UG9BXtqeE3oK/HwUZAcGUkeGYnCOMPjLpoFIWIYbJww6XFob
/84qc5hWjVnA3QUQ1+yKi2n8cT86B4aOstQ8m81nmMzxyxj1wDb5+nJki0P5v1+GX7EWE3Dbim9B
ohSOR6ET7sk9CxgrXvMJopC1HOqJS4NJLC0PMQVFybLNOidEaFcI82rNn4mjUpEZqcFtx87QASlS
5LuaQc6E6Ol5qUMpQ3T7bQnOgdicvuqa8uV758LftCLDEuYzYFD9zWRyZbMFSvNlPAeG+8IBiffI
omsoY4wYmB4svlC2dwUBDzvmWOeRbnqDnRMtjMlbxXQaUELuHtqpdKv/wTG1v4o+mlSq4rF1hLrY
skucZc14jb2d1eeP3eZ4rf2XXw7iaLpZ6Entn3JehXovS7+QI/DvmBkJNv79afKjrQOIYcvfrtek
4XUvbULoOFvGPpjDFS0I/osLHvs/vNZHi0sr8gYU7rcVcZagHHmrUWn0yP3+xyPGazkn9OHTVLd2
7F7ho1g+sJiU9l/kRpRA5s4C+Rz5tHFTt2UDqbPmKWDc7FIqCK3Fo/N45j1JTlzXpgwcNTpsDoqQ
xiqMEaxR9yXD3kvsn8ri6g9b+uBZ8cvUlKMntwY3InsQz88569i9optnfxQGF6Ifm5eY2mmbEbcp
YPPDY7I/oWfqQiF2lBey9sX1O6M2T3H1URh9qG6mNiXGWJI+R1PGfbvkfskzc3tBltN9czp1mO+S
tl3mRGFpMncT9WBfxuukXkks4Fepo4pnj3uLiY9GMMfCbjipO8p6fPr4YIo8OQ1j6QHoXQIkuR7s
2HnZtKjJO7IzuJoRX/fLQ7foWxVRRXfCGsuhZo5qW2TdMAR+YztcfcI+NvyRRzQl0kGKMAmkq9S2
VBsmR/Kqvl8BFvr0zzK3ztLjCPOIYXKzn5QBzNBaGhbQ5jVvOiFkRrAvdq3BLRBVr1dQ4GbsF1+r
nj0JrvKJPz95G88OfyXAeWBHRfW83vRjrIlWbqfLAVTO+q+rRgKDj1rVvXMgpIFkfgJBOSjLS0cJ
4+hjhDwP2NdeIOn6KBrDEWSLC8j08moiILYGgtkyOvkKKkcuN/RMUpUjJ9vBJ7okUx2pj/9aqBzA
sFJpkPd/IuraTJKN93esiTcHdurVVp5V5TR7FkqlSM4da/wtBYJznjRlriWlg8KBtrbRLZpRk6fv
6Ixf2huJMLfDkNRbJPVRG9fK4VewDrfdpFO+Gkh8xjbao0eZZCaPJ7HWlEs7eoVaJ+wDVIQQRiU3
oKZ7nL4umdRyVY9rNc8YN+PdxJi8MJghenCbimfmGJXaulpnlslEfNDQArmSl2GYUU9DrRMKwo75
7t3Zd2N57j51eEYgdKoxih0awrRZ1I1yTfxZ0LLotG0oDY6xaHmfDt0L50GMpdEk1qaRy04qfpsX
M3lgA73qFZXFOrtiil3ryJayGXVnwI/NmU13JxJGpYcCRd6LmRxXgz3aODKWsjLcsyRJna7sAmpQ
APQHLeqPCLEEosGjp6v6aomSjNIbKRUs2hsbqDsJmk7NUlAFbuhoDLUjKNrq/XtpeV4akaTHTLKd
Ywomf3+Y5a5N21x7M08HLMuWl0imQEwnnTsCb4g4n4A1QXCqHLGC/sxDS83NLyep0cHDpXUjIFYp
8rnLi4Au9TNmDj/Si5EMhY4Ts87+hFsRe/6fvR+pctrn3xsS+UPiXEUnPcCoQxm0KlYploovXK6x
WCvqDzLp3oaQgoKUCBr+noZlgM7k1YY4qUJWW8yfHcjE8iMDzRBqnKawwf1CD/vx9XzWWmOWCiFw
xYcZT+2C3RMUoCFsB9K5AZcelVTFJtazukj+dAG1kHMlH5nMeQPqN1sWMvvaz2WpPiVmpa4/36UL
G5GJf7fVG5/1n1e1M563FU0dmONbzIic5x88QfAfSWBaGPaN5aB4FIqakcm215i/My0RjNLFIoEe
7nXQ0PR8dJdMgwpfb19mBAF29bBqWnPMGJrfdW7qbNxa8BToplA3zH9RJp6JrBSQ4se52B/0DVxx
2N4flrnJKOKHEy6XpFwOad/TDAJREBf7QNmoGJx6tW9EJ9CjIaj59EvEmJZH/houO6QBr0Rc1bbW
t1lB4fhwvMhxInwgbuqtZVj/VlcyVM3T7FzDxueIHxI2nIdwKKJSGCeuIzQ45QCzHnl++oRa5jce
mMVU9LZYGrwjKpD/DXSIUD1Vu+2kU0qjK+7ywLwuFfsxZT/qdS1UTb8SVFTXAQrBLErLitCR/tqV
88zi7O/xcLVl2dvQqUVWPS8v9Ux8r64bpTN6vqsvrkL6P6EyT2np0cXAgAf8M0INx/PTNOJr4p5K
NhzrmF27avFuS2GHOQqb6pIKD/ewYlB0uSNkxp3uHmDeMpGoM/kV4xrtrANT2lby/KujgLCWAbb9
sTn+xN9nh++5XN/IG0U0ZwiDbGGVbs0vRFWChIcW+LFqQuTCS0lLDh4GJvdmZRSRsXl7hmMPsCEc
xA4uXN5TLvcZu6OA3S6zjWLCBTpSk9S34pWk3B2p2Q9Of8h96YqL15paZ7KIo8pS08ySs8M0e2ws
s5HQeQYVl0gort677AaCO763F1vEuZabWOWgHKM82+sfRdyI0vmSig0BIK3UpV6w/rkzTDpF9wut
meLUOuAzc09MTtg/mEfbATYNNJmJR+Behgo8lUwyAEm/hezUfsHFnFyhMAOfknQ0GAldxQQGmYW8
/CzFsd+6s/7dYdaCdljf90T4ReAoTatzNLx2ZphWLQNHJjbwQWiBCRqxsn8BpHqzGjWVpcoKWrH9
rYEp7VA00FXuq267dORmc5modNHDyhh1joZkeVg0D6Ihms/HJxIpkgSC2v5QJW3dJkLUZyTTWjTM
pXAh5zhb/P9sQadx+DRZV+DCypymsRArt8Rjkoz2O5pDSwcCC9SsGIS9b0jnGvdnwzXuHdScyc+K
nqqiU85HiKy0ns4vPPlv5zo7k5lBSSH1sjVo0YvuP0OXwpXizg/ypK5tMUSINmfhLM/TtM0jCe5O
T/ARaK/VczqeEhBgXQ5LX+sUy6KT94tkNDPAM+zVlvBPv4O7L5nCIvCBwcFUsKLSEpJw81xLaKqP
04lAjqbMrEO+kTXhmvEE6YMeY6AaJ7VGfG/joSuhJEMJhg8NDsBDDWTwnvhZrkm7Gr6otS5I9wR9
bGhEXsn2RakZn3cl3V2GuXwx8qGZ346rmipUJa8y2pwxMqcAyHwe3mBK9S8F4Zh6QgyH55rACm7V
KMitEuQT0RvSWGnDien5PcvSCDAntLTctRADyyzOzW6GA3Eg+pwG4BArfCO8zbBNUUptV3vuL4QS
LTNLIvJQKHhzAL3Xgtwo14l84BSHARqj2heFAmbWRbCfgobwC7eaTcbNV/c2bQrJ06BpJVEVeyyv
68b9kME6upsJMs2uZKbgsEuDRm9168uCXPXK0ZoKxcrbQPp4ZyZcpKAodPtD2dJC1Tg+QE7AsliN
mv7UA2zpWrY8Gz2cH59kFsvMboLIThNU6SnOF1PAX28mPcHm0BBBJNrBHRGb7udab2ikqAOSAalD
zFY0eMR7Si3xHQ2QCRxjbLWPG0A7rK3StpDTDCOTbkAgFIm483RRjvjLvLU38kHZHIGeh9qSHrAE
MU5VDdPlB4zBUDpOH2J4Xqn0EHKXrP2kVGYhEfiQE0QXIs8UhXsAeC57Gwjs2md8VN2VaOzTjbKg
CNW+NsoPLZvkaF4H5ghm9gfnOhtrHZ41vm51t7yImiKDJslhG4Eeu3oPQr/xvcANbxDHIuRQhsXA
JCYptS5AGBoP0lPMLamzVb0JilZIEkfTa+Hcv6iLVWX0xAniVtrzLwXf4hNnqYiRStLJ6EwgR7vL
NFppIgR5ZO9TU+nYN6ugLrjczu4NxgvdItz83NSfPRx9u2CeieRONKK0WkgKj3RYsYYEe7Mh3HdR
cQaIaLjPj/PpW6rPppLRlBMqnR9uT780PCDnaM5a6KZ5373KYeGx4Se/fqRcNsmyMAmwTjkC7udB
zUGTZjZ6ih/WhxiU64V6753S/d5KXuOYYMge0oXY2CfxiuOlZwCouoyHo+QgKuL0bomEhjrhxmCy
JOQ+5I4fcj0/zsYD/hw1Az/H5LZAvHhtJtpn5S3ocX1VwWL8qVrQGc9HkbRuMSivUZ+emFw/Alqi
cJGFboDTMydggCN6HS1MMInvMNwk81mnjmcXWUVpfMKzr4x48BQrNdXd4h/rapNpH14tyUmVot8L
/gd5SwV5iwu9LNKOn6Qu6L7otsvVYZQOYI2xW/iBNGwFTaJHHfJnVR31P5CXAnDR7j35oQTswQx+
C64KLwg2oipoGq9qJb0fIJVFUQrBL37lQhUZJK8NNZnxJmTqCl6/EmrSOcODYVMK2xLteoL9xOvg
EKNzWzCp1Gq+7C+EFzx7gSJm/BJTi3SUDMj76j2ML4jEImmyS9AArKs17UITFkUfuotG0R99JFnh
CGLOG8LjMzOOk+gGacnZG2Q0uZnj7fPVAtSru9kfp764RATFpAaKGTyovFSn19bDbNbNb0auu9mr
RFHbQFIIeN49Fqstfuf4APXdZ6tdUXJ9O/FBiCfGvQS0+FD4SywVpu57wU3DrImnYbMrz7PJMIHz
BAOU9YviR0MVGQ/rSzzLSH/OnWFBcMb3semnElHhIw1eT+o2/4m4XgbNjC3yS06q6ICmMjQ3qnaz
9noLuJfrRcepWEJRFQRqC9dlSwFMEuY2KNKVn8WZ9welR+b6h8rp8KKf7UOjEe6L8A3bDeky+AY8
7/EvdauyOMzqhDF1/fAMRg2JBkVowd8LXi7paxTzKc9xcQkPC65R23fem6aF1AH45WRPWHlugqY+
aVhNbTQv2Zsf7yyaK0PxFvYUlIOrSI8/1MAW/GnPJNRytfwuDyqgnWHkDfnfn/JJ5ZeQ8LFD/lrC
w5QdG26DvgbWY/OXtjFAw9aD/SR2Uxm01PK6WoEJRglp5rs2jxWpp4xa377Fv8v3VwIptv+44ffY
OHyJj1uPebk6K29ePa58x68pV+oic+LeRm9uEvefLHcBWI52iwtcAVRSz9lKxyO7+5ybziWFHSrZ
lI/EOl8lQ/O5YFN5ZbVInHnonsvPOtdRpGNUzUEccqTN9FnYBzF+kxqMONat+Gw5bVnzH8PcGwDc
BzhO9zmPRxILAGNIdEMEyZKVWH4VV6G5ROyGahJYBxZUvm3kb5llG2KlA+PkcaP/5irDa7X0B3r2
S/YCa23sQiTJAro9svYRkS3N7KonSitdFXv53ZOBjOdIcIYyitBCnhPFsg8vulI+3OHA6AZ3s2jd
ZCt9hIqe07KGmEX9SWzcAizWnc+e/meUvQGAEnKvaqmjsIWD1zzVkISSlLSAL/fkhdZHkc+8bFRT
yY46PbU/78hVHN1BCHXnpwngOJFbCW+PezZTrs9BWhIDQNBxQsu1zSf3h8Br1d+SSht9MIhDIMxX
+xzgvRgHgwcjwbS1CGmp3V1zANYNmI5A1o2cm7iKn8LIfvoq39Po8l1t1nWwNtrQJcTFO/7H5Qq7
AGGgEd8rWlUQ6bzrfKt+fmyjhUj9x33NXwhwle38sNJAXp+JmRhi4WPme2YWFBZykhEOYOR0dZJx
v6Nbvvzw35kaX0gjdVEUqVIpLyZgMrejJUqkm05jjBRAUcWXbWS+Op1iFSA79A0hg2vkub4qTBGJ
ArfGZg5MNzI3zmsJ5+7K0LlYJUkaHhyap70Xk7YsqmlfhH7rkRhKJ5GxpSyFqsshw3TmzBvJxFjJ
UQnBsNP4P5Y+Gb7qXeYXlVphNHhnhFlJ6m4cTXxtwq0OMxBPx26E46r0MEA8HeBEkEuknLyQGijI
LilbxBRhGg0KPMmTjduQWmPpTkp6zGUlyTeeKhKqs1x2lIz/Gu/hrrQBfsuDXBu4PKHP/rUQIGKg
vcgC268f4K8fN3T9IcwjmgHwfK2/MGUsrYQJNVMrUTwlv7PXqWR2lBG5IUCJljm2sYFsD5ZGLB8b
kQqs18CMx2OFSDp77hdvG6BwT9Z23w6Ie5KQLkF2fZiFSttqvlH/eNMYumAdTTFiQ66YET+xPwXG
QMxS/DELWVkXUT62iOgkhNtEAAShBUnOWj/v8FhNhfhylxX+VbD0hcdRrtaAKoFJSsea9mVzJ/EJ
o/7Tf5vT7iKm6AnINoynQlnbREUN+WjRphdwSj7bQjHaxMpRhafE1oXai5vUSDwtAgg7hUfY5Lzu
5AwuPLafqkNupD7GpmjDHPYA7Rv5EDd88hDDZjVdebexUQAtJfnthuNpsU3IWBSdbpLQ89QiPZn7
GWBxkakluODybYcf5rwuVfTms/PmIU6nD3NbHXUf4ximRxyd1Eg9n0yQHqi4Xj1i3m/AnzDRkEoZ
Tx8+4p8qmewVASKmTrbN3iXt60ZyMAsxJyIFBQhIu7Mcig62dkN42Nkb77YvJePCl+5ynuhhP2Zx
45929Wdn6+Pc2VXjeZoGicFZYTdOUgZB7ByInno9ItDSBMWb82L4yF7pxJ/yLj4/xlKILNooO7Z+
yxnyJkF2LB+uiHd33QxdhMn/gXy4PXg2cGd/qf+dDF4s5ODUX1GUMDjbX5SrXrCktp0HFo/A1/1B
Zq8M7pJdi0IxVOZAhtfRJaHqPdwkBEiCftZEYmUuQJ7Wm/kKSQvTizfyNVaGzqouHa1SA7qG5E/G
oPTUXBldGpheCk+bjYlUFFQZlxvJMoBoE3xlcuFPSEbsdoqXDnspdBOzv00wSS4d9tDs1/lRxjWq
vpqxbCdB/EegZJPDxaqlJ6QvSGiwUTP7rGmT+uoighgS+H6b6xc1vcEwaMXlc9Ep88kNMlm6Wz3g
1wou3VmsJNMM+d/pZsWuE+mpDeId3ALEAdgyITiVLlhS1RIGzd5Em3VDnK5LGgoXa6vl377JrxwM
+NYqSJ29A/LzyCI0F/aqfnUwcuxI4inDsTUaef5hdo0s2TGkU7/CElynD9bcXmVHrLAobVo4/ZNr
lYCiPJ1v71mjEbo1UWT/k55hIuto3gErWviWCYnuh7xkeN1hq8bThDzLA2bHjMzyPzJNcbhkx2jg
z5K2fpVOr+VxeAP8MreAFU30OCmc/M6xugylPwer/NL4bcL17pXOYxbF9eODRZez2jO4N85k4lwj
WxIuFDcR4x+dliAmn/ZRzgWlXapHGA9kUdR58TB7pO+ZLfjO7NhsFD5uYi+RXm45a8t7svW2oXhO
FCsPiMiYxIZQfNMyTho8QDr4ccC0ToA6e7CWh5tYTPzap0zKqMwBef/oHoxxhL4iJue9RUmlQdWj
xmLZEdOy/NBSEWeXSBkEOGsxwSRdpg9chxOu8nh/wgwFf64SyKl66C2CLU8vmETOUWA2924VeED3
CJI8JgMFGF1fKez2D/Ofd0DyA8aDCAl0w2tSiKbw2Um6gohQAuf6haOTK+uJZRCi8Dv6hn2CqZT9
pTyPsXrAu4OYxTL5oe5u+5GoE6+AiyHf1aLmHO3dOB2PULn7ivYj5cYf98Mcv3zxz1lKLkSulv7H
BMxYvACQu4wGVPHu27I20obOGgEhXvzRb9LeTqfm2glWNe//rTVEkM20g//eVGewpc7a/44VGWqG
2uhbwB5NNLRY57cZKnXb2u31PdD6+Fvav5uyVClZmPJ+PnyfxWv+VxLLEpeBXR3jLPRkeKz+U+x2
4qCYetOkWXQ75319BgO43mO2xEPcN+o5Nz0pWY3YxTOAjRT/NDyGqm5S4OoTzNYVjQQ0CnZq0X0i
3EFEMcVI0xzevx2CSu+k5Cqt3ETTlUSbmQC2V+WOzP4VvFW7J/xIp9Yi2RbJ85TorolhJseBMiFo
BCiqTSMNhoPSRrH7g7tYg9ZCaP8QgqTEu8lxDVQGLaZ9k/0bpvnwuHn3pYnu+wiAb1UMcTYDHxFD
P4BrkkyMyGKSuoCprRDBrDQdXJj0pV7qJ5I3Irg6/e7yid+SHFSKv+24LKsUTRJIWSJBaHMPcEQ3
VhY9U8EHSQXkdz66JYnwLN3vAAIsAX7rsesv6rrWFg3kDzC4KXLsSc4xUMpSedMsyYWMay7CXZHG
eAwGr6f5Pvv/Qwq41J03bzixQF80CuxLMO5jP7l1oeXupamX7Vjzo2+NY2O41GoLqRP+m3XAbGTA
SdVPRcxogaMGGvTKavmyirSKILx9MVG4EQW5y4UPztJkH5qcnoU5tRvqwmxo+g9zxhvJPXoeUbMw
aqvLrxXlfS0i1oh6MNsGy5Qugc6GscQ3HsEUkD9fjhD9S8oWVxFlqmLSsXUewL8czDmfDJYoKCcB
i0eJQTLz/BHHvwQG+U9o/Pqja/l4WqqkYkWkkB10ISL1q+CtWQKbrHUzz/VoRnf1qZL6L2W+/kh9
jjoRdKm+zUkkrOEr0n2zjFIHN8wuDCUTczwSEGF3dY2VC1uDD3KWttiVtuLdRWXzJ4YiY/i0HqUn
Qg8R3yIfwTCnzITI+1HF5qm/fFVlgJe/hmAdKyhCtUZ0ho3gasLUehEtz+dWlqvoNzPHFfxcvwjw
4pm3M3VroXDk0ALIEIH+j7InUecLa+wzzlhQFvrt7OrlzlZlI/4mzRQDSgafI4w+v3xL3wI3AOM9
p+xT7WXY7+hqwe5iozxqNcbAgxx1kdtQYiRMJm7GcVkxJhDqlqpkm8wTiorQDb/Qw0m9Eq2v5GS+
/yt2UeMjr/rZ8eKW5EqueOG3ziJz6aElpanIy+gU25d+Hq+QuLOsjtwGnxM2Yxsdzq7JOlbKZShI
TY5B/dF88H4cmPmodygHliYQd+ZQiLAmPFdQDUB5rDKOFO2F27EeTMQRLK8MmiT+To+CKUWt+ybi
O7iIFli93qkH7xwNI24TkBI1nh1+qmG5nYNPgSHXN7sO8kB8rJy1dyfvPcmvi1v3GlHz0P/k19du
BsyeC88n7VdZgpFzHxamS0S5yoMAtig+PuReLyiVQQisFeiF5Yzg4tAf+iSNpthhn6a9ELMmyUe7
cMicsXYiZv6u/UPZkE0NKsCla+9kjBNL1qKorQSFjlH9Y9kKWRthlGBy5bczIEH9iYsKcVO9QHdk
CILZMwM/F2RuedSrYomBiPQEr0SqkgXTcQ1WfKV8pXS7dZoQY1cUSo8XoRrfKwhW4t4pG/l3e5gs
3O1mpp2NZwLHdnh07AAS+Hl5OhfBM6Bqg6Q9z7i63rJGPyiPl6sacU9DNk99aiDQdlQKdFZlNSrv
hEaa3xkanx5Vz0ie+S2AOy3sUIKr3Mw6C/iBYxMyA9L6YtBUzxK7wtiVXLcZHPf1o2D5Rdv6mG1w
FQg05Jwu1ZP5W1zVnGyNfDmRFRB8E0IjtBQrJEzNdmlb+MEmbDhOQ4jTqaTzu0b/xZoQqMKTAWIM
4OQEC3Q8BNAggKnq5IWs7PlpAQE2vZ7ndfddYI9+ZFwB7Nl3G7bm2w9XDEGeSOzgOejyrq4CVIcy
zgVcIrNbYzmcyNMIjCBKGZh01BglsIpnydaA7rKlk3yQeKwUXMcwFyHha2473FUnm5BjLh01MPqv
w5bPxmX9Ma508jNb4Arl8bgOul5a9ZHIuGwAJnp6X+vsogH334YAC+Zd5C3vQtofyyVY0NbUabok
/d9WLDxyHkKXUjwHfgnrUopKdOTX7cI3t+0ERDYcO7PHZ3vIxyTB1DgM9zrP7FDWQRRL+bLt7uaO
9Oc+jbM7a0zMSq+et00hmhAoIrityn12MNrGMHBITFXXu7dFINN8FOjO0CorC6Fl8mMzPOnmuY8W
La2DoRpUTxKEJFV4RYA646J3PNaf5HEUPxdQG686zrPnjJTMjIIeOdcNtkH7AE48gvaKqvsnNJvr
RgCuLNBCwOBSxZMTuAfzCljHBbA16AdqsRTGQZLdy7EqG59L1AbqktJs3SoB7SW8x/KeBmEoNAYN
tSEt2oERDyb9a88zEpctcB8Hn9HTc+tJbi/O7JbJCmWXGc0coCOwsDwsmn9BS1Rf0YBOA5bviA8G
EjeJbpwhflr9JytQ6gwI+aa0pLg1CvncPlsxYP4mjgHra3Hxkc8fJCoPkdP98cYWhZ6zbKAG2Kep
TGrvCjkF/IzwZtOimpTm6fQstuiN4hVSGDm8vHaEwHmFjP4N1ITCjDu3g31rtY859SGMG/GBtWR7
Uzizhxm/MKLZdSnwsufPkihU41tbu/n6eUKfVtxtiaRBKsWNzbH3hQcgb2GI3G0KPUNEnSLIscCq
oY+T27MvCxN5gTAohFBjcVchWfy4qCgTAE74/BNSLTEazu7YqOqOcSfZKy3bQvOHCjLfcApH2T4Y
dSRk8ddY3pRSt59yHqiysfAjzwC2pq6iLvBID2RBIAYj+noh61cyOCj0iA2rbJyU8Tziwnh/tWwN
SELiAmyhO0q5HaQDzyV1YRrgePiE0ygfDn9Zo+Gg3TcDPq1XVnF13yydx75Nyegj7mDALtQqY/N7
cZcqy/tVKRWONTPanUa4pI2ZB0X07ZUgLDIV8/m0Y/o43PtsZEY/roVFUI5HoPU+Vx051ZVvTX5j
kTVzXsPW8uLtDCsuxD+w3+6dfsQVpS4wCO7BJ5EAdT+1ZanVxr7iHUK01pKc7/jAEt7kKX0BxV6k
T3tBXdmYclo7Mhtjhp3CjFEDiazIC/13kEW6Q79jDwklA263T1UQ/cWTiaPlRIe9f9ED23NvzYto
F+YUugyjoW8Lrq2dRHpHGYFA04ME5fspL5FjjrvDIBjP4XCy9shkPIWEP7/C0XNoNLZNmvORHMLh
uCODVarQz4Gpglg2ZqnQvuN5T/YedbsMRdC7GjCU2e82krxFSRP3dC8gVs/eKHWV5T1KnRp+Q0BV
lNUzhq5g2Fr2vO/zbf8GN/9tq7LCFVkzwkDrXXj4J7TIEJBm+u4N351GA/6xetO8SnlHf0/ghR2W
u8Y871PpgvO5V+mLOKplu507GRkLvT3PwzK0dr/+fY/Dxj9uPsxRfjGJIxV0YZ1la3aa1Gw3dufz
Nt787o4EThipGHhYkj0JrUUgqZ91j/3Z1wkt8s6fVOqRrYHJ9+mLMA8b5bd9iEBDJUiS5cN6j4L1
h9YmJmDxuBfWLJwhNwuWxmqItqPxPYhlA0Zxlptq/N7PxaJ0lkEDqwveLGfjfHi/fc3kph8t+unx
dDSibuZJTxZ+ikYk6NMNGRwEXKxjJAWGe4Mr89dwD59Zj/kLxsHeWq0Emi9voEoBhNAyhMwolJMt
j9Xd5lKZ0rT8T0yvVeLxZD6itrZv8e3589LZ7uJGd0qGW9e6fl0w5CelnERiHEL4T94CR2f4ehu8
dqjv1w194gMwilo5eJS8zF+7A1bxbRQECLI8kdJC+VT+Z53OZWMMELEddzoppo8wfFdHpWuQiu+V
9zzpz7I4tcCfwVLbgScKhwKjNcahMFeOtG1mmqqpSXQgduZjqf1bJloccl2jeDJ5nKfoM+y7mdxY
RYPbq/1z9ebT9/tKVygnuP74SAAQVlQZDBhGGrJLwv0GgicQ9fzbLQI+pqbegkOc9rAjwbZrq/XR
uqQQIPHylB25NdfK1IICPLoAKhRCLdmCU7U9dD54iwbtZO81RVGQkfLb6S/U9B9JYycDJP4nDuoV
3k/AUqE6SIZ8eFI+zYNqIELJOCT1uzy2lsviS9ImSH0vo3GMkp9PJTfFECGsP/iQuOva1cy7OGaP
jp1I1sbxUiHzSJkqcNJfJO5ESDZijQPQWLMD+l/7OhAsafz4VTGbv2FGWaQm92tHid10bcCTOUjn
YkYOl4Ky4cx7bbfiz1NPfc3dgH6jAi7cShqJ8EYFgZCPHch9qui67+32qXSJuTCibjjIB5VouEGy
XY5vMXLEN1EzkzJfBeVk0ze8LFgwsd9NBgbRCVqlESZcDvBjcs7DRUV5+4Ih5P7GNqSYanFx3NCR
AyaytlWxOBsLnf0g8eOoLpbuQh5MYT1QOmRcWswSwg1xovDQoVFrDDkuJNs1FTU300dIaNVqJTx3
lSF1Vr0ruSgi3AD5g14tfXAdyy8ouaZvv7DXRUTdd3z17HfbE3hFcePsc2HFZemgVQ3TDZI833B+
LPZ40cLNQOFKons2vkoqTwO7qlLZ30W7TEkZ4sbOBdE298QZp8C/92SzZx6VBOF0m3DBbkXJK2p+
Kks8Yznkxc6JXY8+2irzW8Ct52NYl4JRkZNFrTkRJ2ufQnhbkAhftAuPwgcpmvQjFRzrp4rllRow
RNT8A1oJ8GSR5lp4F31qSODdSWxwhyjxqH3Rr6Eo9o6GbKSNBN6vonQk1bF6UALG1wMvhpuVb7yX
NRpjQjvpXe/hADXpvfeHQwvknbCapwbo6Y8l3t6HTK9wh184Vvy/pq5wkupaMItbaRKaoOMXSEIa
9tkwYEfBwNNstNjZjzt+W1SEbKZUSxROUUGGebeh7oQe0ZsHWd90HsP9xm+GQ5Ju7Mh4xHS29tKj
v4hDCmRcrtfDu0Edi5/VWN7PkYZ9d533W7b7IAjYI/MUcTaw4CeWMSDseZIs5aWCiJ5viK4IVHqk
WA6g/jkUSyim5wCOMviogUjzmw+9HZAa6kLMjy+K3hgGsPSr/BD1MksHZ8mqFAkIEhbt9wZGSKU1
Uj9op96llJe5uio1tuGHXsadiSTMcNqgktXs9ZXw8cv+0F52nHtcIDnj+VvtnJMFBIh7p9IjYsih
5Mb5+cu0yTXKV/3eiMjvq/A2veqvAGpOqNDzOSKrknlqCfi61R0NNOA+DDLzmNco00X2nvB+wLD+
8OJmG9oAbc7FSu0csibTgqnj6u7NqiSPLhdKysO74Sb+NaYBQK1RwCeJsDrFtWlVghfubym7W2gs
cWAwWluHMqoPAXSj+KfPBJrk7EmyfPcXaUXhCG+zs/SbeEQhp9OpAeQYuoHRuf9zjZiquSaoloqP
GU+UEQo7WIoGwG0N5wO/f0dOenOeLy4UfF5ifcMI21fsJSndL67uS8Q3dsk5mUtlz/sUd8Pww4uo
VQM5Zdonr9rqDyini8+jUC4OxTqGAANMGjQPP0R9vKcFvOKEnxhX5ysYSdkYV28wt6Quufomkof0
8Dg4AjGiF+OGczcaqgLDeQ5ewpxnp8kaGFxQsjYgbln03JC6w17MORE2FLkhY4YZMLoNO+jPGOtr
C+8UmjiGOKUAThampDUtU9dEDsQEUjNYKMR9upqR26C06Bve6caYOObgAK2517fEY5SpMdOb7jkl
FrKt64GXydgMjDuI68mLYiPhY2lQml4LUN0lS4IydqXZ/HggXZo4rscTSAXSkyZcb7DbjmHgmvDQ
mBeCMJLhlDE6Xs+WOuhXzUG91aoW5uGH5+JrG+p6IWCJvyQjs3lENRfgY8MeDAPHNCKkyZE2g/ta
Glh7FH03RKVgsS9STb377IaLLqONEGNgMaEeD+/ufd+bs7lrQiSjxHJAnQjfUhJuAG0ZK3sqdhb+
Nkyoim7hl2xNyARAQI6gtbSuYWQKOvvH8/TO+EwwGee9yLYBjXO7n/Xz8wl5in/UzItrkfaL8JY9
5apRtBeBMnPJSsV+KLPQQvdj1uOoabWHqhxeepoqmOfLPq0LNGUu32r8TJV7IfXZLr0p06O+vbXH
80gxgLOHnAq/MzdMM7OcBJvCgWdZVQV1NxeiV9uefyjeYKewlgxhL++QYG30g9sG0LE/la6ghtOx
ilLzWptLTD0J//JGM+o6pYE4p1yV2zLwirkPqddGqHuI8bdyVKiMz+o5bYJKEcRfgOaWNGxbHuXt
kw/FoP1YzJyMY4Xsslw6XbmntxEsB4N6YjE/6VjUgMEVk5cWR7gy1Ff0/rTgSk/WL09Qq7mhMWku
9orColpclDF8kO2r0cjyNveDq5o5cB9SPmDxOO611v3b7jeVACZa/Aw7b15jtf2t3Odxn8xpmC8h
pT5ewihsTwDZQKxDMFPlz1ZtWAwcWQ32sYX5LphFA+tgM9XF22HWZHkZl/F1Txua3fP7xZ0jjb3d
UssedRE72YhGMD/buB6kWo5ersTHG7U0WKdY06XbcI5VP+XGjINVThlDVNRB8ZJOoW1DH0JUfoCb
0dBJXuf5kG30He/4viX+irgF3kJCGTDxHqvfPgpjDALEdn0PqU011wKxeVGKXLJqzN2kXIk9BMst
J48t780RNbZ/T+bqosV9srSffwS3pl1jrObnMCKXHt6vCfacULGr+uar6iDE7YrNVojQXUH8e1vA
xPXBbLDsaEvWx6ykUzgouE+MfzOdp8q4jpkbMSN6uiuvmBeqlscNTwko2M7ZgoLZzxoBSMcKG2hU
A0Uq9GHGdbrOFB6dbuYG1HR8rYFRbPNwXsT+En+ZbPrD6ieNztNnOdhkKBeLi1AAEIhmWOYqkTGT
KEuFHIY7v3N1Z6V2qQjU61F4ueS4jjDO0XCgVfIrtXZ8xztyOOz4HEQCZmRoEhAnF9NRPGwb+/UP
COnj16yn+FTWrdGdCWKfMEdwkJgnXy/dXl98W6V3F5AIeBbtpKNv4f/0K6TV4mRS58ori34nCr4Z
43nDack8LMmf/C3jP/X5W1hi+3qbRCSnDPrCiFMZvQ9Pxgnt0jR8Ea1GRy182mq3YcFZcIlwQ+Y9
J/PyxPdVfD7c4ufCP08IpqakVYvkQfsE5SO3abHHYg7GJJyRH2fzmKUAtjO/nuM0ky/2Km0j2LMc
TEb5sGq3sk547RtD1zydfh0ovgjLsbg+xbiHOcg4ydoMO0k1lYx7jFmcjTjpXNpVSJzjfA7wgFdX
UrC8SIh0J07NGgJ2UA/ejjFQhdJCo1obxx5tQHeUy3zDn21wwP1AewS//NX+RUHUkNCJmwQBMV3Y
osLs+f6aWidVoMhfWr+PXM1dtUMFDTnffZT+D8aSwyjIilGukCpWHmSVPo8DqXQ6ujEJI5PyHyO7
YPiIb7sgUFuntjUaHT9Vxe8zQpzKgruGWpiRPeqyVOZPbUYYv6Gmx3wRQTF9HWAdaEn30GVJl+RI
WJjhKMnzAnt22CCp8nreLPB9YsIAjxBe7OEDQWNC+vayk+jSX7UHOKeKWzxQ7ufNJV0f9NhtQ7w6
3UcsJgacEroqHtQphG9yptS1/v8aLKzn71slpDXbWCYkRXSibQz/6zuwIvvR56B+QDiDXgVS7JXX
t/w9c6UHJNMT2wz94azTR+MTfRglGJkyF53Qpidgl9tfBJIbtSpoSIWvteDmkzNWXZXPP6b5w6YQ
FTkTpH5r5d+FVndsfexL3KSlfJLKTPlwaR0Q9S8UG/CHXBY5eGeCtK/5ZiA8v9JveiN+ICKMnjxw
l9ylvFbhJCLTFYzl/lrEhARqcjoFG+EmoFNLfa9LMX2IDI1k137/0KjFdzqDwqM8192w7i7c8xhf
IqDJDcOrMLGuMYCVe+hyxjTAl7aahiB9Ck9+N2/Qo62YCAmwF+06YT0estNSWns/xMxyqo50/Z0K
w2stGPpWOve3/ZRfwCOCJvL3WBvpiKBS3Ktz3lfWwfqGf0QIty0W3KFQw+VsSlmljknbwDmgzqPa
z2LaJfLTEK5WJA6EBjnNvMEkdNTSU6CqXhy+BxWj5k8BvR/3kpBh4b7DTAeIOd2MdzQPGcQaFBqU
rR0lEwG/38j9KSKAIoYmF/bAsNGlC4ROUawz0SzrdsXmIYoSKkbEdQvylaL+sT3NbWrFlT0WX0Wx
NmQVpp2MRiOqIdRWrmAw+Y3nBMYBk7rYjpF/PIBNAnuuUqXPg9WRaJ/t4VBuR0twt0dRgjkJ0w/l
3DVTvANAF7ureNXCAaZ5F4PYWsEVMEFyjdhct/CS6Izy10MPPSb6znyCSlK3OzFwivfnBxyqvp63
S8Z7ltrVWpHGLcv27O2XLjdQuOd/NpCnrWnBGd1mtYXHmwN74u5AtJzacYLDUz75bR09PjN3xkFK
fJfLbFd7guQ7rBtwPOjZzQfJdrLK1xsF7SuVDUPARREXREVU4Rtlo2ALP3VOewi0nTFwJp9bF66H
9zu+hzYqjOIYBpBLzeIjLjug/55Q7UyAhJQqjbminEw07iRWdeDUPNJrHGrn7JgE/Ruyz7MeRhtp
xxNHZNccTNuZqLxTM2zmwnbh21eZiWbOqqw8Xat05NJWe/N0MlIU2WkLhznPo9nWd8UpTqZWnRga
amTQ0CZHPhQAeP6cN8g7TwYAGNoqMda2f1WQU/RhMLjJ+4WXFzVjdRCxmXpGUPg+YZj+TU+6XTGZ
8Gz9Dbi2QHIVmmaDgiQKwgY+UlF+Dq7J2EqxZAOk5axOlqwZ2qLDrPfN26is/TrFggBkokuZoUg5
4weWFdmiB0RYEFOpDk8+uuYGFrTc0F2pjx3RWqOiWjssOuLDuH5rk8h5sD2A/RwBwR8ODVKkNH0j
t6c/TphUOA7Igi1Pl6Z7U5FpTJdyy0Kop9ccoSx1kdCa4kJmEUsNR8AxJWIGHEpreKKhDntZ2kxf
CSXyUkS5kPvNjNcz6ZCqORXdzWA+BmSVOy1amrJAVbDUBH0F9g43VfGgUgpk0CbqVILx4+FveC70
4ZpaSKadFAJAgwfXM0HrXfpxPCzQX52D8vF1fLsrWYjdfFJe4Doy7lP12kTeQoE8/WjIoiGpamUi
PQyDyzeAxWqZbkdNGIw1uWZrfev+dObXPdxm69p4OEhEw6widK7Z3gBcp0CDKpS/g7AjzEAVIWpD
v8PWNTCAlG5eGMilVklgBWkVG8Kz7CJMDgEJfYK4puJklyBcbx9KEkHqa1uGVw0xY7kM2I+3ZYTz
Bn2Py8HXnaEW6nlVTUPxeel23ED3DkTmx4MtTgcOzEaBq43ha8XMeMj84aueVDTfGGSY6VbLf50V
oblMOi5F2Jsq5v9t4rbTOq1GWCuWsKVcySbtrNDUTX0xFfApLCLXPhJ2KmzZ3k5iM7GbGsfnrEsW
knKVbKky4TqKHi29H2RoG0HO57OgyKv4jrVdi4AaIc4JXLy4QVzmOPVJARj1qwkZNL/7X4EL4BcG
UdToUEWS3HwLr5skirsgDBGayyhnh0xGBW7mWV9o+D0FjFbHew39RGWUohHNnIPl9JeiPFq5j1rv
Rroq6DiEwVUPOoqn+SjogVR3NK815R6LrHab4mMY5hv1sCOA8D34E+0TRPzQYFXtvEXRV1IVOLUL
ezyDmzBTvI39BNn2WEoECTMwAmyFAn8FENkLRETgXy66dZIKvT/loovqnRfoiRpVYTLVoSHsgl2/
u6eaJMRoMOr7AhhdJbpkv8aBwN7IQuOHV3rfJMsbF8F7/SJCKFRYrZiqpqMXXhay6wtP8f4GdYF+
acqMCaDVLMh3fdmvvkU6gESZesjm9OgxvE21rFSz2uPUWtZNILTI4uHmj4mtSnBr7bCBJcFy2XJ4
0fuJaTU2YjClM1BSS3F7AzuN/+lpoCP9OBzLl0RYMSX7Ie9qT62EljtTiHubbwJJpSevtng5woxt
X1wTvQa22l3VVjbJ2TPaC/NQfBxoPzAGL237zYKQQaEWLC6cpNEb5hsUPTqdaaBI+DMpAH8LTcbk
QeBSz8WUrCfdopScOVyDpTXbg8G5L6/nQFNzC0lWN8cKH7jlcAXYc1Q3eGPL2HBrdMXuhCUyWsyw
G83Ir1ZzNOqyzdokFjZmpxSk0yNtLXKNu19oDwX7hKa8Rowcojf/CWSjIyaAr7z6i9v2IQY7GmZg
VT748XPecSqUN3hQ4IHTDh5c56zW/H89/xUu/MxNde4hT4Z6k9a6ojdnf1nHs1VJZ8KP3hOJxiNW
oUntqunbh7Bvbd2tRgn/xIIW2uD3QFH8NT5BmW80ValEhEpBc+RVj5GqrQqC79M1F6aVrrcW7Xdh
BrvYeZOZN0yx7cZda3pqQ8f4ccAshKpaUwPEnzmRBNuGqJK0sdUwsnNV9BfaH5Ahko650tNHpTFp
2ulVTbx0DFlHiNa8newY1/xu9z9guwT+f/llZLq/Ou8Vcp+2boWzK78GCUgvBMLEZH5eEEsVG59z
DVsYLUJxxtsA43hSDh2mtWrLFuR4CbzODD77MmDlXjkRmAhqIdEuFGch6xz+0jwTq0EwZNILoPDy
JxpbMalhLAY5AswyIo97Zrp/J644BphcewE8N1a2k7vbMA9z2rphqee0xjG77WK6KBc1UpzLSwcF
Af3LE3ZtD79SB31JTx9CQOlegrmywdh5DyjP5zNQlC9sYFJxsLmR8N+6YIqs1xscs4oDfipE401t
giExz7K1H9D6xA6WSTkDDhbjmQU7t8cGI7txUy1MED4YSE4IfnmAx7//dPLvNxevMtAw7dlipkH2
9RTX+RxljW2G0sQMgjg9NJkKf+w9qeNY5wNSrHXvmX2/9QeLiAHCnoJmcfUcSmx99JCXGqC8gdGg
C0h4TcKHNJNS59Q6MLiSPwflrdHqA2PdPPAyZFsNk6+2/rpDaePInSTTLY6Z+o4vGsGgW7/FosGX
Byc2IE4jXcArDZiodTLB7cy4yyq4U7riQZYH2v5PjkYo0Jx984605m4JO8hJX1MqhWYEct54k5wm
EnRrfp0oe+CSYxDkKe7Fb1UjnrS1021uwnxRDFdFOa/0eLkGFM/V53CHKeNHRZ2OzeMLZXluPpae
fZAwXSgNQza+9yQ26MMQswSwepJSf+wISaGSviwZENh7qr7OArAvKAQO0apxKAEOA6qDT1Wasqn5
yy4LlyS+rC7VPMUXyC70PJlVf2DDVA98KcFdp4rYApMK5E19SoVbyiKiUXjtX9TjG2zT7ATfxF58
n6NnsjM+YooyLo7Qew0SlI3oRDcrgQaGTfTq5WovVpJAkDQsgi3J7CGVc7aGiQEf+h0pli5evFIs
Z615LtNZoQZeRepJ2H6pc0kBVgGdkfc3WPO17GyzlB5J8USu9JQaijQ51o4EGCi018sAf3VV0QtC
Hx+YfTRZqHTs5oNoDdfbENm3YzhBUzJQAsR3z/SGI4Vxhp7Zyqz/FM4zCInSWDDD5mO3LhXOpi+H
Vy7J2vgyLgTitmKgU6ymUgVR8Mc5/tLE23TJSLBGhyudhyF6c8mCFRWBZ5MjYBs2JgloWynxKhl7
YWFa5XgmIx6KhbnwV3p0BpXO1MCQ4MjCPu8QtYqDtLW9aMi9WDPkzfN6V29Ukt0DiKDUyKLfe7ZT
Bs13VXO1PgqCaijqKBjjPFt3e4cC7Eci6cq/Xsbk4C4Bi0FgDo0dGal7KLWqNizA+AHTlj23f+mX
8Ja4RuecMYhAdZaUfyToSHcP5cdRenikyLAIQ035NE+N2voZiaHpfRHeGpy+/Pqn3LaafFWat4RM
toFNzjvh7cdI2fpi1su11/+rYhNiANnGt7GHzVS/TXzmekNxNpl5Yfi1QJzsh7lmo9yBIn1N1b5a
bj/vKlNJI22osRmEeBLL23xnPc/d8y+/jZyh/8z+q7/C/0bVUdjQjkBBoKrTiqttYzy7nv9pBNkO
C2TxHpziYMXt4TinEv3fLAziruMWq80dfbSrhcGVxvNCzS/32Ju3ksx7ZWE5bvnojncZFjQM+V1u
G9uaSkKBI8DFYNzwXcdm7gYQODeCCNwHkipazK9xXROPVvJzfyEmzHVyy26aVvfG0Tbnxc4QsJ87
nzTEppp5DbKe2Ep3OlIKW5VUOAqIhzOdo+rKbANbGB85vNvuK1L8gm6oDDxmOTyC0pAFj9ihBXct
+YnTwTP46RDrEgfbRcom4SZzsKXkfV3H5Df8PDHb5aQCakMLa1/94FjQqSO9H+nJC3DjItIqsEhy
EA7qSRVSiXdsJRZ6raX6O2ok65qZUtJGzM/4TaJsl9UCBjUzums9ahAyHPeuZHv6NEhZ5NobUK28
odc7lsBtZGK1jqUl6irvkvGSLWiEEJ3hFUo3iOhQc0YSZGSX/m/jExWvsKn7imriKewbi/cSSWt5
nJtquE5QBF3ALwF2F0bX7JFYZGQ1doBu+DqqdwzRHt/iRLjoIr3JfsnteSvzD98WD+f8O5k1CzQ7
EI/z+uNar6kipmZKR7Jubt8l9ncIu/W6JQomKzXTeqJKdXmoqM+ehVWqm1Mw+cATI9GaLEm1GYS5
eO9ecfH8FI/4mdAapYA2ROlWjF6vb+7iXktSqna87V8q35trljl49FdqCceOBNsP+H8QnKPdlRjj
5zgtKwGJe0+wCJ1SHsEt7hUR/Q4OkwZVlQWjB71xmswt0cMk5pIwF7s7Bq5lpkDKg5djQxfNfgMH
Z76MgLgmzcLvOHjCQu8or8NluAKNFtlDuxtUH7Gkl7FKar8fYP1mNcdWoHQoIS7LKB2skPbpqFvA
IQ0cdytNp2dLfuM8TcLEu5m4aINwWNjJD0NZ2KcboixhJYQ6ghf0OKEzGQOkdLFzbEnrCamXWT1G
KbZOT++OtQvnfnp16Ho5ZNLqxc/Hput22vrMnjMhIarW64YH9zsrqxS+EMMrnY0FSnYkh+1xjBke
OmCUHb2jK+XbGBiyEkZujQdVNBrKOL818EW5KOfC8thuXqfkTZO+lvFNQRLHgD3vbhFprxF7vPQG
cBqxMh73hEgug4bZRTua8rE6h4je75Nwozwi6xra3rebC7FUMMawJO6kXf/zsAkaYv1nXUZOW55o
N6OmUc9bq0Jx41rrzytiSqxVgIpwevI7FkCwmuEglPwYST6PGiIg18HdeAYin4vfAJLrDFs+uz1a
T2igY8LV7k6q1LvoepYcI15Mn7857lcUXBHfr3K8xSJc5k5+b3l1xXd0v6RcYStLdwnzzxMgeXaL
/HZqre64SX8/HxvD9IKbyID7tT+AIBoBMKlRThasg6fyKudZ8owJQ/iI8R9RUI1hdAfqtphXckg7
QUtMZMV5auk/zAryIiNIsi68ILajLP4eGcfNhrS+++TvUE0YqXmftSPWaoTPVZKBjpbG4vtpN75e
m2V/RHQhoD8cnpmoqNVtOtDuZx9B65I6Lr9Y3+ih86OdN8rKGmdAojFwJ/AfVgIJ8p2ZA3SZuZ5C
5bmKWrqkAzak1dSi1mhJ9e6O3UG8GuccjtUK2EdrhXW7QA8cwohj7hNfSPo+O5izAHKNHIOXl22z
74UuYhrA0Ki/PTjuctwSxKACworjICrPxP3+fQNEc2c7r+eUXdTJHLoDpaEngKumHAczptO65i5G
F2pZjG6g1Si+ENafTS2H/uL7IqY59Td9Fti/DOeReAyWy8Przc2SAwGsLEqP/8N+B5jK9pjOA3Q9
nGTsiDQHhrRs/7NCUUV1calbiqy9MuFvRH0/dAhGpR5U490SHoKF1cjLTAs5b6cCgiJlwl18tMF1
1/Dn+8TJTv6A9boTyKkdSW1sOMjWrPIktiEE+2BITaJvrCQHXDeGPdjokG2NBKt3TyznrF6M6O3a
Om2Yebw/e6/971r4DZ16sPcOPG7Q8CeQ+PaM9IP9DwCC0l2w1V1bvjpk9vinl1Jfv32hg07MgjiT
zcV4RJSfW6zpuRHPwCBxOVJaNJ1qAj5JGyGustLopeoA6AEppMQfBbbv5JdFgnxocuslqplt8bMx
Tvhb42NnS25yXsiEAdiX07pVjcmjf2IA+06E/YxG3LQ7rjl/sOJoIPiGCetKPqJRKOgAJTEMKz5M
BvRX5QhxQWK2OgcWQ1pKbPxJzZk90eFy6aRNeFr7g2N0f8htN+IWhfcknHDF7iB8yULC7jJzMWZs
m/1IQvdDRiNpx+Q6rWrUn74HHYS+4Hp+7kd+6gpT+gziZgXFD7Q/nRcDa4LAXnRd6CdZ2RqyRI0S
//p+T0XVbZqgj4w44b3KNu4VY7D0uauxBB+XRQugx1jOYyAPFpETEBEnbzoMu9Kc9cPovWk0n4py
dA8Txwbp0DbNF8Hd4htwE/NOicKzf6N38mph9STGeR07qDNhisEtBE9FXtpewTQPUvCOvL2HOgyh
pflaIznDY5MARS5GIqfRAhI2E6X/pIHGEdbRxYImG+oeCjcB1k+G5SOaTn03kp3veP8T7dpsAixH
0nBSybegy54aP+RnTLeK7K0QEOqe3xY+RmiM7H7j0XZbTYdohEy+cpqiCHUWojS5rKJ1jM5i4V2L
tKIOCrPLTPQgBtLzo97TU7t6AOPFrDYQhPxRHyvjqiYG1eZjIiLCpkpuUfcPpqrxZh6I2Y3vgtvN
3gdP9xC5DZK0l3oy7z2B8gxD18KEVoybIsIySfg/zKIzawhRTFX9TW8voy3/IYgF1eUbtx/KXZf8
NuUYv8fgLTAvOhvrjhqebNA7howjN6N/cp0V1mZ9XwOcliW+G28T+vO4aRsFBVa8DfhGAp78lLpf
W2yzrpy0IBoiJDvCYvAtxePb0+9hPoHhIxyBHQA4K2CD7Pu8g9AfDYEvM+yPUa+EB6bycDv2VxsU
Cwy7fNsLhL9WdG5iqnQe3q66lNK9wzrsIX4bu5xRhHBi8x9VA9Id2ns7cKB5JSJvOx/LXFT5FNcT
4ThAhY7pWXyk2LFRUBfCHiPFIQdCpWJbpCu/CGtTrKVTIczxUAid9SrIi/pZ+vG8X9r00ZZtkfy5
mNYoC2Eum0Qqsdq8K+NphmhDZNZuYTs7dlwnEbfxutg47VOwfdyLpaOexQ3aPtZvw/dKl6NDNwgP
yLouzB3ZFn9lejOQVNrV7SeWL+3qhZgt0Nq/Ex0oCmFaZHVn2gO6KLAtKQupfOAzIeNtapmcvIwE
m2gDVnbCDB9i6x2ap9Vm7vMC3dY3WL3CFIXFT7HiSc5w6PoaaDIJF3uZZSGTvJY1lFmFrCBpnKpw
oVfs1NxyNFsru5vRzPyHjWT3mNaLoL8PBcSEcVhZhVOvtcDj3pqmBRpiTulKbCScDkmg3ND0Uiv/
Qr8kBcZRZI1WjqxJYL//pGxeLSutaIv/Bx5PEYPcKqmFm81L2xHzMpNkM8VnZqnOIOhAGNuxyyq9
07yMPhjevhbglBVM/rebC9IouTGCl5f61BW9hLZr/EQJAyexW39A02sCrycraKR07HL+LZDjiwv0
a8uX1/pIQM9XkCUH13vFyPD277MNyIT3G8ftPUGQ10/F6VSEauNg7LMmuHzD04ygJpMyaM6BY/Tv
VyBPU9ogW0muJJnafT5kZCrtiKtPRg9rVEnKj7fdJMkiVA7VqPLvnQ08EYfRurtGGObiOA5Mp2T7
/+vDczQoBy0j8EbW4dd1JblNqcwQnw5kskozkZH22OWKt/Rooz4F1aUDmR7XItuiKTOdpGfbhI9Q
bdZsSj9bh3EJAgUkf0/kCKhT7RCY3bjkgwX5PeW/yluDuWKfOVrBUuYBe8NaZheckV8fktR2eZS0
Ht5I6UsfYz0Co7DMUxQB+YicpPJUJ2c8HDQFNVkcJhzz0B1yheVTSl41TJF2qWS8Ox0rLh1U+0ew
35g6iN1+wt1xIVr7Rxu6/X+LlVjPNr3RjWz34dsmdIB6X9mhOhuEmhhZdoIg/rjWU1/zPJbcq44+
uDhuvOg0cNzmtfPAHCb+62tfs5qUFI/V3FHv1Jk62yRUifVFTufxUUM7wVlfhXv9Lyv7/atffeAd
FrOmoBNZpoH7Eb0/aJ8ZVshOufS6IR/YztCjbqj0WqC/ckk5E26yyE1wCpz3sM1lNpqsKw4+hNAW
bXdoaOqg3Q1LgPcIsKzoPf2JfZatG6MrHqrQExFJjPBi0gm47zjTtDxd4PWSgW/lsbufuRDmozDL
acUTWOnpcvYoJZuy4yVQ6BsW1b9qfdZ4FdzIo71oPlnjKlvL84JlGrOHpCZEBHKcPMR3Af264hhr
JL3Qv68f8BprPFEXsSqZdMGlY9ZZfpP3BK8hoG9mPtS4jRv3jtg3Px785u2uOJzErurihqixQZXn
FWzxodXA5TSgE2ZLUEH9o7L/5aGm16ypQyAf1oxwzK3KV7LTHHT1KqCBPuib20FkxiaYtB0lkcv9
ZRI8UdtiFfSY9PGrSiLbB/jj37Rouz+3K9ZF9zaBChn1N5C8E2Yn2wjQ45evDcL+CXcEh8I7jbgp
ttEQFQvOpDFm7GFXCzKHlPmMC7MiF0O7CeVRNKyjwd3Xrm6CmbKdLR6fcDTFalBmppNNY36t4pNh
JZ3LihSxkNmRe6ETv6uimqx4agaND1G9aPe34xm5KlYOvNAxKfS5cpV6sPNHqsM4oGkpqs8O4hXz
b84ffUzdRXq7QHuUAsYURx0MbvlRSkRwrn0rGys74AYuDE225kLqTwgzG22oLpJ4vK43b7qFxSsI
07jcoERjEe3ENQHxv/IG5ae68Qe53gnj55c0jve+sIkbCrKzPSoKNtcrZjlVaM+oq13yBaiA9P1I
87I1FCijzeWHbOsIMovjknu995M5SLerPepbBTFB493G8+51eqb2f4tIx/RqcUhc4ozj/XVZbvyP
kmGVwwHGqRY5GMqc5mGzCkU23iYmOwIfou06SX4LOtkUyI0OArh9yQ1ngzYZovTtYS7G75iFmDFk
PA3tWe+GHDmld5ax6njbYj483wugNxPqJ2aatbY3R2STwUxvM9V+nzlCXkv6Wh3AIUy7fvYuJFsy
7nVgOap1QMrzSmPlob64/pxJLOqj4Xc+L6pm08qzl6/MFI8YDCPO+3i82si+4c00NbnNWd0KSGxO
7/nG9lww3JiIkuUbRXgREe5TIZ8ivwEg63IOeWFyhWYrXMOZ1bRQO3p+6BEnMJHdwl6yL3ktf7Kp
Yaa09fsQn1o+HJV1SU0BDkYgenjHAFtOxbYyQ+NTDouc4GH2MQJb/eSVISTKvnsyfl115S0H6rNa
zkcdWtgP025r2So5eGd8+qV5s3PHVTZpKf8rjYiPs7HHN8PrU3JA1fM69Iv70dFJYoxNr5idqYrg
LnZA4leEJTh62vKWMqA4BjCCbyygST1rQgJ0HN2GwONegzBNFzPpxqjfV6jovfrKSL0IKwv1kmY9
ieHoEMS1o8XHWiuo1/p2RcC4QaE/ZcBMaP7x6dA9gYI+VAF3dNrqpe9AfqXU2BfDBqXeQlVo70jl
WNZFlcyLQ7rYZ7IVCRgnKDt08eefea1Aa83V/35nGsiL/wXt8VDcTwW5lCtc/rgkY7CY9osIchQO
+F0nrkVDyh8RtCJui2wsqQWCwtWZO4onpZ4PQD0HfCl+b5lr7prBlJpAsgkSBey3Mw16fqi0ONNG
QFxx4/MQBrlGU1l1Sa6qg/a9bHdQ58by7WcMVvaDc2Gh2xjGbAfEpNFpZVfKZtFA5KBhm1c9oVpg
ZEGrytvF6iSmAxQcYXrD6SrT8AGIYAj3Vuw0gKaM4EfGYDt6Vs4QUztF4UG7AK4W4CzQ7meXVzSH
WlIiAap6+b45Vu/kZH1H0DAf3anFDIDfVFG9894vWZ6xYDd0nlKw3Yq2T2NSJlKLRtw0yY5zHeNp
zrX2ED3tJH6K5zv+6dLpI2QvEOkMD7AvitmszvHnjiiomU4v4eUocp+EweLr39tWAdDi1+7ABfta
vMdB08Ttplwu+1XfLf7iNAlhGpxuG9oqKHZkR5Zph1KqoTBJEJuBn0xqN7YcxyqxGMWKyX46v6Hl
yxm4hymvWL6mtg1VzktTllAnoO4b6G7S65sz5lp7iCUXE8z7aixGjM1Rg8n6t42Mj9vzpqCHlM/o
6NqIhK8rPmdCzpAfEl+FbRj4P6Crz0PKhzv8Ej+MANlsA8sFZFcVMDMwqOQJvFiwqah1iJXXD1rQ
rOsHkAT7DIceGTBNdWkSsva17BAYa0T7/9+uoy4XxppfuetdYmcNlat8ByM6HLNdH2LPeb6MmkIk
ZWhXEUGHzz84vKBxQL8QecZCCts5NnDFH2RIgtRary5YpMC7oJbwvop3wbAtj1G0B9pRyjYz5ish
k/2eSTd3PXPRaLSeGeMlOEzjB6JmPQtMTRNXjt+RO6FoFP0W6cYSGSmSMTghEZcV+gJS2wYZesA+
WtcYNwtVJALtGx6l2l5jq3OPdSNnILOBjRbW/WC2yQBgL8LvPJrckFLZlMPhsDb8eyXeob01lXCm
CY+8ElPSRrLoSBDxXqJvuhtnoiarG+Qw4AMkF76utX22bHJGpl8BKOvON4hqiaSQzMXvMw07Ql8D
Ueml7xd+ksGfqsUctIziohdiQsSsUQM1bQ5xhjH15FDVKRHUeftH2BLQ+7xBZCJiWfO53zFBxobi
lHAuBTKGIs0zAfyGxIRRYlQgN5CSJq+6+bMZysX7cyopw5NgjujWMpW25X0B4c2aKQoqX33DNhp4
bP+FFcG9FUxvcDJfoSfpjMNxDWCLK6hN066NU5uCxkhMclZgEACXdLHflAmO2iJhDF7Nkg7neIwz
Zja5qbivrSWpH4FfJAOKZBMYCLGp+NIqCYZX4o4CB37sIIN0bPJtXLMP9zeipQpbWCgXv3KB7C0O
mVIwy2LMUtoFKzt1a3wTNd7YUznQH6ODHcMQxoeQp+H0e9mkQ6/81DZSYMxYAPe8SGaxvcphAwiQ
Oer7pGHKn/2z4k5CVpJtNiIidJggRcKTOU+h84HT9RTpZnDOL79EoB1OQyjjn/Ev6Z4Fbf+3EMvw
8Y7Kh1mr8+32FhAzshRnl2x5B5Vpf7oH71ADO+RtSx8THpLcI6aCWXl2hX9Tm6sAVXi4c0XqBsHp
/bofap1Li+P/J+cdlAbVjBh+rRiVRbSW2Ur1mfr1pFxQlQmzQfd3XMNAtjSHse7zuIICHMEnoCOo
7O6RKiHKJ78qRscXT7gJjDDeiOjQcidSv0jcO/9U/jf9expt8CzNBh+NP6uDilVY5GzjZ07TMKZ9
82qUnPixN7Qo0QlLTpzb22qLdJKCyudILoxxrLTHEN9z5QW0CENAInZWzklEYvaZ8zlGTlBfOa2f
i0lJNoVdiAnD3e3mFzWMpEPKuPhO3OrtAEKbIvc+fA1D6F6x0EQsfJwKYN/Iangitd3EMNaFD+eE
r17npvSay3RdGvQeGxRkRnV032Q+oo6iJEyHkrAPnRa4lYstiAHh4NuYjfR2XFdkYfmNS9jzjqUN
d395O9KRd+yuH2/oqktBJeLq+SzbkpF2whIqFFArw0FYYREtBWMXKOIUa+sQp0gyBqYqqq74PL+n
XxGP+llwbulCvrcJ3vLJtjkyCCb4m63XBHSlLPb0UoA/o4xYdvapryEeFg0u7/h4vR/MQd+8ufsz
HxKYdV355PoLX1xiWMrb/1qoCm72EJTgOCgx2SufAC/nBM63ZLJrU0hsDnhDtUmvExkayng3fVqt
EH5SGBqN9+p2aWWF1VyYZWuziN8IA5uR2Fzsfzikk3cvLILWD1L02U088LOtnUM9WiaIrGaC8P/J
KbuDjJ8GeW73E4K7Bo0i72r/GGi/gDAR6rc1lXsl+xAFjLBrhWnqa/dqy2qralPlyZNp1Jfonc+0
I8tbZTtdZRC1SmBZR1XhJX7bV1XL38ppdS3ivfQsFcKQMDtN93ZPmxI+01hqRqHkHIOfIt1aJ7cV
pD+KumjyemghDGiBejOg9I+ZQ0Df0B4at36Ju6+DTFhWuNRfAImsrqBzGHvpNp1PIrIX+U3D5y4j
3nPM0i6z6XwDpS+Yotuuo5W9A5I+rrMFoWaRPszTwJ21Nkyb+jE8SkJMglrlf74tnVJJWdKU9xus
Ci9WlbXfejlLWm4MmtX9moF6gon/vFaSSkLUPr5T5VYadvO5IDzRHZCOG5Go55gejnUfS8SCnNxt
yJobXYNfZ6xh7vjOz+FOUr7Gj/HSlFICAPWFO2pR2Ef2s453wQy/vKBqJUv6/1ep8df+oRFaOeI9
17aO7UnhsZ/q1TIhCOQCOe0ZSshdcPXb8it/NrZJpqE0nWw5IZVztsxOMNf0kHXPBc92tv/lRnB2
bv7lo6ojDP/uAmN970RtyBCybQ+cfLaE0thash6eJkBYVeOJQIhn9DExZ78/VfdTXoS1RJ0EHS5Z
vSj36oYq4LdVYyBYLXw0dRJKPAJAX8CcF9U2PILKXPI02hxfHKcn6QO7GAMeIaEtiJv9Pgg3dsk/
so7npXB82yW8XaG8GC5T8A/vcTvf3YudM/MfYP1hWOR6eLSeC7K4r+ydeJxBPKKOIRs4/2w6244V
jD58qzGBfwv9jbq8zEcBYC4ZHLpLE+6REkFGPT6/tZNjpPvkSwx4G+p2F49VU5R3xblYByEWknHt
Yjl9RE0/2/h8fgjZWpDvfpfQEOqCmESbJcawmLpxOwO9roOxB6VXnLHBFZHjD+eeTcTORu1y/p2o
7l0/viRDKMZ8tGflhoo66ngFRZ4Tc9MPL94Zw9xpxJFSc3K73wN+UI1XY8SwnQ1wr2qcs0/xYzpl
XKPIYhYZT6noxqB/g/1kWdXO8xxDb9UCN5G8+qVivPzNV6Th5AKqmDXiCmY0iDqdSujBbquZKgHl
nfAWnBdULvTs3s0Spj5bv7FxMjIpNsiPVnW8t0/81VXadpZqQIvpAWJAOnsz0eq5IjYLKgsFjzx1
uRPBWSPEVqRjKnguTwVMAAohDwOCLRhxDVpYiGUfzeGS/S8z+h4f/vJziGNkFAWyYH6LWR4hI7tn
0OyBsJPqiNl67l/9jn7iq2SqPJgNAYrgDnGe5fjNwQVsMUZq6QZK5FKk1lCRnABbDsY81Credrez
2iudS73oUrwmTfZV8/CSQaFnnfHuCuI7e8n/QmftNn4+lT8vxfJ2PfYVMBKJwFwOKJIVpC+36YVC
Mm376xw1m+NECu1jyHEdjuNcbvjzVhHoJ4akWpRB6pDYDyfNlrW7yIPzUObMmfLrjTCI0zj6heQE
Rvs8BAKI+//e+c2ny5eVAyI3P3+/vyTT2hPvo8XeVTvqjYPpmySZyF0BOMqxPhgvQLhwTP4pzIlQ
m71ktQ3vJMWGeq0lrtR8Gw5qCFQmDKYE2uIHeG0MB9o+ycxNSl8WPInMsnwvrvfR48YQGn3Y9EZG
NMzqppo/ZGilycOlsZZW9acQypAy5wBDc/+VxxtR0k8GbG+jRIH5loHiXoc/09hKbhU+ybQ284R3
bFoLuzLmKbZlB9YMujcmALnCcaaQtNkMaicCWuksy7Ewvb4IQB8xwhY9udp78E6DNxjpvw2/9tt6
BRhjskysS3u81SxjFDPYc91z648COU6fX44nw4CvA4q6q40avqMFOz88D6kS/KhKlBMVfRNuCCT9
eWo4jmzfKdvYtO9fGD7FiAOLvov7M31z2C3J9otH4yjNPx+6mgKE0+r5d3XI2BO45+rHxgs7sUGY
awwILF4ilrBKRUN8s3h9hicxAWe81PNZ+DGCsbjB0fhvJYSdfaiXvMJCGPNOYC6Px+QmYZF4Dsjb
5hM8ta53nAQQ7tj0dY/o+DxEOa73Dc8vt9nvcBzIC6nZ+kFQiCvy/MyofgFij4ada8OvyMLt6xHS
Fz+9ilGPVaWpKzMACUDqrADs+OmtE94SE7yehWuoAgU8ZO7bYyb4bJ+3bd7dDTlE4CPyHmqiHt9x
ZRBCAFFUSuNFXYUp6kA2NbUcgbCMPGF2NkWqm52w3lHN8d6BcFB3D8eHVM+arZd/qxdFhNwmBQil
V13pg6ojB2Wss1WJbGvgR1NU1OdVOkJa7BbiEY3celXmnzs2iB5fD75ERiYHoxNRBcYOqdGJAWuQ
hHm21mvIfXxLolazHMksMo2eKb1T6tej8vTrT6xWPG67BVTAxXOeUUwdT/0MtMVOCxCDwUfd5/qd
7/e5mfSb8pDTNHheXb6Vl/Kq/Ry962JeUnLR7uyzpcyXHXWOjQZ48suFw129LJ9gc3dAPs1/B3xW
2tLS5R198K239t+bjzaR4Khat3jpy5q5BUc8xff99LAyOA9BAGo0eitgze01DBPqqvMWMIzHCaqI
b57lCF5lO0+ggINnaKKqdeq87kL42/OKMWMbVVu0GmaBdUcqZGhoxbgwS8l6xfhB7PsfyNEBcQKQ
YiQPwbTX87dBS1V167VKJQZKR8igO8Lh35R6tPkpSUjcTnobUUmxDwURK8yondODICgPnH2nkw08
t5hyIKL2dH4PyNLtLnMBqjc1ZLSEBnT+MRdop5jFj4DZ0YXroehNsMw4q6VCg646kvH6n70u8jfH
etZqQ9Ma95Bbn4MyDIsLX7iwPXKFXjNwl9T7WYqJEHSRJytYWprcNFkHDwfKQxmcAUZelmT2/sLL
Ypa7tjEWWbuIxrzojN6Bi9lB9w2zW3+78FHd+pD/ictNko02yTuvSekiaSvRce4pwDgjwiINxlZ6
ETZ+svOFWnjisYNg1w58Wa5eESk1+fcrPsOJ5i1L7/HMS0XQOIHvZj5oj95wGSxNWXtk7Rcc2pkK
ytEIEg+KRsaKPZtgpRoOMLKSaM2Z9e8W35xSN96HI+6u07p9c/aZlWv2zgUttJj0R/9ercdbDRlS
0QDApLxv8Xkm+le7aEbHAhARTsUh5iF68rmTt2uhaZRc9h1Ce87AM+Am4IKL0xmeXjl9o1iuuGEx
QZ1yDIJocG9geBU09XzYJAdxobZyuopF+b1DGpaXW8pRlpm07ElD398uGEu3JetWSXdR3wFhls/D
hEfPKgJD8DFx/RXYFsAbyz4Bt82XRaYK2Z/V5JUJsSpcmb8yx5AY8Y1w3muzEdT5gnENvdW38N2c
utP1Pygtfo1dAjVNY753mUtjLfg/GBZl5f48MW3mpfkcRuds5YreZlkyLTD5H8BOm2CE3ICaEzZQ
/Wns+Bkr1PpxJTN5fGLfG+avHR+ixXD1A/9861yGBV6v6cGmmEGFbrmVHaerYEAYzBpW/u0C4ihD
KYqO87DQqkJs7em2Zm60SlkoVbUkuckXDuWtdmdRcfjRWr24W5f3UbmoZk64RsuzgWebcmYyFic7
jsrDcD3zUFtyK+Uh/v95+aFzY4sW49mZVQoSIPW568iLxZ2RgGb/6q2tZmddSLozXNq3h8tn/Jyl
rX51HzyWPzIv3EuqaVEKvN0ryTfqbNU4x4bL2tAyoCednG0SocGbi+rwpv21QXqTOT3xdZLBQCaS
EnfsjRQUn0APveRpX+rnN0WpdfAjKUo7jzeiqfwA7oRkGh5dzoKZ6G724B7roW97BBIyqGA5VQMM
o6pI3tUT2V6DMQccOW2FLi3MdWWJg3nakAWfhv1ngn4vQu4nqBbdoCxcnEmwfwUK1ocvhotnePy5
TJxsbKrkzELTQPweY3GZsTYifP7/7e42156AS18mz9RsY3VvdD8TnngPBTtxciNnBCFhcF3u7D2S
i7Gi2f+UXwPq7xfVGJuJhyV/R0EnETBxPuSbO8BCoGh+oL116MESInRiUukK37Q3Af3l8m1y+LIa
rfQh4yDdZDJ12aEOpH/wgd1jjDOQUJDUJfpCyaqCHUUQcn0v5tWM3ckcYhwba+g3VJe2+QtbsGMv
9DGsPWdwGab+Pp5gJJbIIFGIO0gL8FXLyxe0Ls6ZEt+oMtl6KuqveZUUeUAQz4NX3QmfesrG5WJ0
2qLaQjebQHNb5PYsjv9T3TbVuvlzkMYgPyF1YeNxSDqsSYwbxjHj7/NvRrtcOWOScGPx7HKJ9yEj
hO6yVPksE+GjQx+lhPD3STp3B3WtYwk9f6D/f7OmQkAW1jst8yQ7pVTX0LPRoJB8/qzHUjl+jXc2
uCQTtbILhAsYXMTyV4TZPpTtKDH2KOutKZmitienBYbdGCG35aLyzXH/IOJu2/1id9aTJvIbQGpK
9zOwUlnhmZZEEILWR8cVgQQRuTxH9bBD2j2jNNUOWkpU22jFO3HR1t05OjE8oL4pVwFOI38EXZzV
frIVF0W89Ep5jiFZ0v3zxICgYk9poGE3CHa+2mbGsQpD3W5x5Yz+S9o9nbyIHym1OCHNudNw8XRh
TDbjyRaZPb1yg3gZFEqjX2wiFsCjPBhyfM7rb1lVs63Ndh8h1R3Ms4Fk858GBN6N2WIgHdLmV4qz
LmtzEGZMebVIBceYgVYkKUnScCNfiSnlGeo/bNjRDoRlL8zqH7vv25n0CLYE/pLPzQHkqJdnGqMB
lxK2RWYuaLLhDkuSTDEJQT7Nm3H7Xp9z7vKTp1X0zHBk5hI+Sr93NThD0xZ8pOlp1ipoyPOqadzb
rQzottU6j14no/Arqw+AQRwRA8gI75KJA4jQ9ShWLT6nxO8VDAjbsjrIarePcPhBfCx9uEd8WLzB
UL+8uZYqfLnCOEOAUwRfbkLd5yYWCIAA8I3tP6lVtSJln39aArc0IuF2JNOPFjvW65VjrcgG8XsW
M20w4f8vsjdehj3E0k59zPIVSErlxu2LD5Nai0ku8Sc5S4zezHOVsl5AjZxzcOnySe1JRhMQzmqi
DaEiVX+tbLXsyC1Zh5gnQUHjBtXXJT1kAKhz5QomSGJeWsxVfL9WRHuaOfyoi4xknmtvukAmWQPi
9JR8JeunNftQq17YFyB/AthbX+OdBkztTZH79mCwdr6YIIQCPvdA9lDShaw4TCxRnuATzMh/KNpp
xUzTnGWW0h0JKBBaqn6FAy70MaheQ5Hh/dCNTokSUT+/C9Q8QhKbPOKGgBppPsgY5ap5tYVwmEua
ZdkJAuq3+kjruUBgJFWNTAXNk3r64hvIsfuCCd+0yHLJkm+75TAxAvva2DcrLV215NVJsUcXCzd+
nNYC5NIVymezzgLAVBt/bv7Xl1MO3Q0O59TJLW9qBf/tm72iahj5/aC81Z9STpGvnNy7dhWPOyp0
R7lBuh5JG/0BsLcHK8ethu5AAifeYhHlzwZjLuxIdV6i3JlQIGMbg5OAGEATxu/jOPsWqz6kOd+W
6sJi12Buq+cka8pX0DZ8ObJ5qEzJdPPJ6B9jnfJJkGX++sCO1vJKTLhRa/KcSpBjs7mSCA/gSQLW
6Q2sr935hdKRk8ctZ+hnQjJDPz+nuBYB3jOw2QFjjiKHQw8RgKOx/KQQQdDcIvxY/4nSshjbppEx
3qbBBE4g17PvVzz+iMPztF/z3mGFGN+6ELqdWPMclX5W2pkCh6DlcNyXDbz9r8hkHZm2OUymVrOE
Ey3y1vpApmZlD7mNbcze1PdX7Xb33piO5zY63BZCh9ayvh6OYGd357QUIaqcGM5N2rZlhK3MelZm
WrQRwP9A2Ppu8mDZaPjoZTlVFb6VmT2BD7xJ7hJuYGnrakJ2f+brQeFxW8RrGG9lTzP+gyHxWA6U
mO9/IVjAALZ2FhZmwAamNEsoY8fTACjlJYBBYwx1eVaL7Z75bLLFVrJv6BUd3D+/D7yGKRUNn0iq
esKFmjve08IJpGVGwvh/e9jTp//rJCTNrRZlM4wYtKsj8NR6+qVOI7di/uQ4hVIxRsa8mSpTClEt
br+XUTJ+3ReWJldHYXzVcld4uw1dBOb56vy2bm0siuZRAKgSEJY2RIAwkEH3v5keV4gByo7dE65Y
7d/IyBkOWg0MbHcog/AC2aGqiygod0dyLmXQ5l+3GzEGY1l/Zn6ZsfTU9ujEcLOtB5XFnocJPNtr
+gUGl2rxTyx2+A1uZwSB1daqcMVMDgeubD4Bva1pSplIXiS4T65VZPIRdRGyGKdCyM5SerG5vzdO
vWLJ1mHinFs3BWRsKe9IXgNJ+Mz1qx6TJj+7yDSZ934lW0rnlCZaLiZPoQIG10nksvy/KnEQMMFT
CmGf5bJ6yHObnOxUYlhMhq5RzVvnsQWdif8dmf5lrU6gB3VU5Tc+FLFg9LAHcKSWrBISMbBwRiEk
feYk+sOfFDORjc3rY7FDIb0KeLXWRtuOLTIwSoSnV37KgHiE6tiL3IUDBnFPEKbg/q6LXmKRuL49
8R8SVZJ0dVY+EpOUsIi8DdxOgdPVW5Aom1/UqbL9pxFyTmqZ5p4P10Cv/FFGSkGtkYMZxB3Ue5xv
8H/L0Dn5F+UODcZnY9alnslIxy0SsOvt9ShVtqpO3PeBAMnuDf2XDI+f5YvrBGlLyMuKlPJhAysN
vfpsYlOIbozSafvIES8TAMmWnFqJJClhlLd6LosbChqI+U/wRjTJAmF1ly/VUkXdNTk5o6QaoVR0
Gky+wqAu/Gel4KXrTKNLzG1vdOkW/8AtAPGdZ0dYEoXP2kGiekfTYahAlPQhKOcZTuys9u4Q5y1/
XNbB0LF+LEeK/8jlM4QkW2h2AyyAhj2o7ZEeWKEQv+vht5B0zgFlpocMafvyupyfGE7KcEpVMuIN
gwr+sb0t1GZ++zWKJVqgn7jxSjB05QRw7RizGJk2V5v1UhjlQTTXmtgsW9NVDxaQKuxHi4QdII+J
rRHsYrGWERkA543QD6gEVICXH32aUzdAWCTnQvzGdEYNNC35OEK7sbEnwNkSaLaUdvEZiMNnAp/l
Yyc8df4Aws7Fbp9v/UtAb/+ayKIZEXUjdCBXN7y067LvtHmkvaeQW8CWKXCx+4ysBJb//LFIxyLp
BLgYJLuwm+FN0LHIwIat+Ts5pRK/jAIz9v+NiXXaIWth0uGOMjSPaIHb8OnSLLFoif73/PQsN+sI
uLeDKxc7uzkKDfwpu4/4tVDtKkQv59oNPFVCmfqwMYcrt3hj4xi67cCAwnDoWuthj40RakejgZN+
X/SdD2F7SXxJh3zQyQbB7GDNlx6g0Kk+EwCnD9ffi/0l4sQYzeouloSc1DGwqnaFixFLmyxD2CKs
J6mYTywxxqg98o03rJpGi04qiqLrraH66uNKxqUZdBffMjtICmyWz2QZk/kRbzWFsWX/fqtLT+Jw
uLWgz6RyFIJH/jb2axPHG32eueAzl5GA81llF+ut8PefDw7VG1p0lKHfMV5lSWcu9/WHhuy2lS5W
W6ws+6Z28F6wdFEtp/Au2a6zSnwRQ4qtwCLQOgU7+j1zhzFM8qgGxwYPcwF6Pzyeg8vkLw+NKRHY
3PK88woBdhtQ/3TQWPRCdLAaZ0EjwSjIV8Cp7uVrLGYRgmzELXAl+FWDwg4RBcO7IlWxErn8rE6x
xL6dHyosELz/VszgvoBpAp8cVUq3JVP2nQ9EuAnckwZe3urFhmp+5aS+5qtVugZhzRK0TsgVe+PB
Rcdqvv/cvGmvKjkbTPkGLOYyn36sPdzHExzCKYkfXv2AMDPmyM0dS6zuGjJ33ze+1hEx7q4cPwCT
eR8+Gd4Dk7Qn/UegbJ9knwds7yN8d23adO3YGPvAU8ELowoiBVKf3qbJL1FIK7wEPryTsYTRQjqK
9uM/Ke8peQn/1OIMc4t1RY6VXkTDt1TbGMo3QAyVov5uoy4Zp+CE+B9lGr82b4WKQvTp8tXLbS3v
mEhaVHXgazgNPgr8xxmJNVya3alaeEKRcZoD9cuOl1Qjdc2Hz3ng8rmoti1owym1BXZr87d8IK8d
V8So84TL3d5LH+mbIbLkes4UIy3kdbp6Glzhl5qvMPAKchxAS/7dMgupfYuLSErZSGzpWUCGElWI
ZPAxrxnteA0nN0T6GQfobTa5KqdrIC4Mb6DoRVUng5i53dz2NOBTnWxrKGSw74dkMI7Fqw9zaft1
Fq7LS+ElGHfYj1AQAoJM0T34ZxYjulHpOhqPKYtCk98khh00UXDyxJAfrzR1BfWYsWZJW4G9spky
RQG/OvQrPCf6ADHqDhYLZtov4lA5qWC740ofplXIDTNuXYjdIvvSnZodb+HzA4dJEc2QYs4uEawI
0wQodrUk6mPOmti5qkg9Pe92Kvnr80bteIK2Fg3HCFTwK1YhlV7m+tzMjIPmWEceqWrzNTwMyYBS
8MsnD4HAsa9mKWrxkv8h9nOVW4ZhjGOVdZu0wEwqfIVZarFBZ6Fs16YyPNM43zzwCRZ6C36ixWOk
ZuUXt8bYvQK72jTouZFViEnlpCWBmMKVvX06NWmxIKW/nlJHyoMj19k+ha5SOrDCCEarIw9NCE0/
5lyDyFU4OiIHjGreqdq1mPRS6aPKKwgU9tsGVR8gwKoxeXIMKn0GwmNH64benprHSJr6uKi53wTw
fe7pCQE/sM0LIxEF1xvJtuGK8QjPElvyWbhyFxgR3qtkODHWWoOGo+P+dPTyZfLRi1qERxvKR4yV
y5QVGRIuB7Uuqovgjows/U5JHA4PjxIcgxiL2UAXLZa+GCsI3mijS1l21V12Wjiv+gUGzGRvO1YN
GTutXJDnWJ2MlDlQ32pO32qpWoemX3xNvj4CD4EHjYUHSfn+ys4PUUV128B60cGaqkvTiTBNNavU
ObQDuyMiFCfBxyh0sd2xbg5+BDeWSstCXUqdE6xUJ+6QkLm6Fve7wx1vGC4PXgnXtLMr3DLZuUVq
0zOghuEYBl+0SYnO+INLpRHOO2TBb7grUYP9cTWqkVNCI6D8I+hLn+UjD/XfQhI/eBT9KsoXwlTQ
0NordKtefPJ6z8P7gQuRhpLJwiIFQ+8DXpn9ABKHpi9YkqerGHRDhN0F8wvB1on6nbW72IuSywRm
tfMyl49N1m8eh4q/PPyaX4Cr6NZCTbg02GKKtA1x/Y4kT7JJLL1S+MYGFxhWlmgMBTcf1dMtRnx8
moB9YavyeoMNc6b8sc5buwh3bXCy56iDonTqgGyc5RcKk+SA8Byf7j+zqW64k+kl7W3/7TOPpwBF
Spt1wTT2s2RTe9AL+AbJ5jfjDlLRMS9rcw328EavoGs//S+traSBtDZkxr9lLJz0Mve2gBjbWfnR
KiL1b4rLHAt6KWJCU13je3rfHOt5qZ7ZR2TErx/A2QrCCGPUOC8d8OuddujmrQm4xGeY8ZzUW6+4
/5Nw7m6I7na2IjySoCMFNTfzSWdF5n/bCaDLwM2lFofdC89cFWMFAlSBo3+PvD2ubVDwLtbkcxOD
5Tp6B1Ak89xPULw2aKeFevIBJPgmKSrG7pcmwhUbsbZNahbF6BazRAd95kmnQShufPmTu2PucbzR
mpfjV7rvv3xPmeuemd2GHmeNJPCgSoI2x7qYPWlNCndLItzPW5zxMdHoFpdy17BbatQNLrffVAse
fHYRg6UOqm7XcXtvbPPDMBI9DwWc2Tgx45PP7m50m/Ya22slKqTOTVg3dUJ/pgcdrHlcGGZLlwvN
ZkeXLguciJ+jxayIfreOWiiCc5MF/NJz8wZKpJWdNJV3yjhyl7ShuecduN1Ylb0xaLJSP+YBweJ+
zeAxSr03I1OXxJXr+tM6j+XqtjOrZvHlFa6xqtHbnTKZh3ZMNBHapPNKm/UcOn2+xrxM9TroB+L8
LSj/aukncPWuotgpRN48igC6/3nSMl7OgyjXhoZz2Lc7rAUnANLKEjfqoLMW5/gPd6o2xLmqIkcA
zRhtKNDPtbcTgtUB/El9331qhzXM5p7gd+cEQUejQOo1Dql0uMs+PtsDgIjFVXb0w4i2FStVQO+q
ygXweMAR3s9L3rAKh6orgbIJORRa5UbVP7tXlcw0lY1emYF7YtHv8XxBkE14Ux5XwFPDm7EU51Sl
P6v4PkKxGor7wFQE141kIwi2gHLLdTnLKWFc6gDRhLJ8bnq3JMSGukx7vY8WmP/6lK/dBkIibB6D
zZU4xI/mw0kObV3ELCSm9gsGBC7zfptsA0RqbR7984Q4dIiJF2/co24F3Y3z8JX54e61mu5G7BJj
DDd2vvSPwbV5wReY1yFBPQzn7dpQxjoOeCbu8NIA9uUTOXBLv8ItLhlPGoJZZSz9EWqO3Wp3I9VJ
BLvK59N0/XxLtxZwX3iuGoYzh/rIg1yjg4+V3TzNB7GEK+LiHG35AQaf8q6fahUT7ahaVK2t+AT2
MevMQosxoeQ1WmkUDnRnFuo+lBf0uVUH/cuCkKKexcR639CxQ7RQYC/v4FINu7YEwVIC6KVCxW0k
6RTnno4r4yZPG01RIGdNHyGQDnelsV4+dZ2erzPNHEsOn7xtyhC+59r70amOQ8HNF65lHPlxX+Gp
a6yIoKtWHXJPMGVwB+nk9m2L/HZm+RwsIWtSth8KYgBqsrvOgYHdarNOco1mwGmZ/CnMXRBpNYrY
7Hk/GLwcqmZ3goW80rn0tytfjIx1b7Eih445CBmNzX3WDW3e57NiM9DemGw91NH7OJ/r+BPIDuUo
pEmFEgRBnf3vL8ITo4VYhfKASve3JFfvrQ16Vj8gT7lcLMs27XiY5FTQy3jSIpkQsP1F3aHbSEj8
w6lm/XQil73x7/J96o/5whlY8FLEt8lvFQeqFnSJJC0zMcGCbrCT66vnzq5LNTnNIIwZYE8UmeQ7
CK5sZGK3x1978UcY2YcTYQxVgyRb7kwcZaIgyQRmiTc6+wi4f2epMVZczk9H4P4qbhIi16lBv8Rz
PItnC05Nm266wJdpIJNaPJLPkwuDSWzOwckATXTao3DtplyQo7rgADuqYrSB8PQ8nGIJNl/Mu1XK
btVnhO0SFpCItj9/RKHwF0j7nn29x4WoT5+YDDgypyjzBDvDfCiqWw29q/ZFMv17IEl/xwAy8umN
luJ4093T3Vqy/c7Y5OW+EFgJ1ON+oehlm+SEIqcN4J9EufxF+S6B42VpKFqYv8n0gzAcl4N9yOW1
dH4m2/SoIOosX0/EcL0obvVOOtmRIpCwZSCZdJ2F1o3ZcZnf1FBnTKtRCCdihZVWqJvmIuwovWVP
ryJwZ8Rweq/vuAhYylH8aqee8MBiq7dJClhs2k75drb5xwDJzv4gdpzQ3OAjW6t8EvGKcY+nPzRr
nHY0Bkbt+iCSvS9FT8BwAVhQ2ctdLSDFzuUvf9UR826o6COF72JTU5YMDh08SQAOM7tkM3PTma1L
dWPb4EhAs8H7qC8uSdfWGL5NIrc+0y8nfQ5TONNVkscD3reNSj+q8MUMQk8DNFCHGEZXAG3UCqof
SXf6kIu73p/JSHGyfLIPyeArSSk0LjchRlZWL9wwgVudnvPMcx/vSuCFP+wNMTfbpzqjmCI7qfNo
dkokwKiW0qMco+NQU108JRaijXPHXfi3q7IbO9psOA3Hbsr0JSO0neRJhFmXWp1AP+0ojn3JF1JJ
MDlCuGtH3sVbKm4RgQQynyFEB9Nu98AScSNr4RB3rMLpOkYXdXEbpErnK46ffRPPHA4otmvjvM1Y
hbJwdfOb7EBVDjqAJP+Bm1EfUlP9YVfjYA/ZhjNqv1lD2XtGHWXC27aQCrVml/0rbQ3GhKuVU69K
y6X0l6VgZnwX4q+8kzbHLMYTPVk7L9lxzr/QQbPC7JEE9P9kdPa25VCSiR3tGThmVbGDTWWtA0Hq
qccODh1udSBIcZf0Fs0D6PkhwCdD2IQ4Sn6uwxW3sA3dmk5REEMUeenFFB9vFdWeT9FzmWikBck/
o4sPqCr5kKFvDfPpJEq2odc1GwEPIe31Dy46pIyFGCpeuEJroKsbU495NZxrdPPFV/JOqPlQ8B0O
O1BOkyKjiSlsJsF6kS5UcEfQmknoiMBLjulTII3kBuOxrZju/Ep07ET0JA+oQ44/tDP5dUHyl9AC
gCjHiiv41y94/3N9cEYQDoZoJqzBQd3GMmsTvzyI3jnX6oHlqTny3DRGZQv5gHqSiXpI2rEsgj7s
RYTkT/8FE5cFr+YWYwCuXy/e2c3IlcqZT1b8OMwxxEK+59OEXsJ8Qv5Pxqr/PW3sgrmdqJGUddIL
5sTEiEkTJ7WUu10vywqBUxDlLcIaYASTg8AAdu0Xb080CeB66RtSjOAJNcjS2XDuuXy9VdzDlcql
NbxSTkX5QLtoXIzPTiiB18IQ7gS2hXhNH+G5vy+zGYBjbMZ0hp+lwPMgegqx6x/Jc43iWunlYsqn
rPZIFD+3krkDGSSOd8e5OsD+SKdzVBL56ZOga4Axk08yUcW5PcndJoaa7YTSLfnuCT9Zdjug6Upa
nTurCxvAWQQYBNfd7oHF3HSmILMOCSC83fsv6W3G/y5Vz7ifgDdiZXaJvtoUrUplhM0BflhS4+G+
uJj2+pwMwm8t0qsqovBBoibzHyx/YTmLzU9xWKgAQKK9HrL5okJ74gE+9amRrrQynusNEQcFb3tK
abBMMWJVnn9OnaA20UdsGQn7r87oSxLn1D8G/KxXXssXQkas+JiPFVGctqHI/DsNOqXuR/UE3RFu
qLJk9su9UPOlOcleWA92tgrFO2KGezjyQbqrYIS44nQ6+D1ah2rWwM4uaXRiRS6ZiPsVNzyB33J9
NUch/9ZA8ziLv2Gn9CUGsG3ydxPBC1zt/uqMiqDnXwGoeMPflbZcQp0O9YBX0mn6WGP+apUKUDAI
To9w6YUSHokQDzwUeW5UZoArzQbou6M9JlHdBPU45IrtkSuUKdzOKlpJfuskyIf/2Ye3Uyti8NUT
mqZ2xy+ypZaXSVXaOdCmd123ITQ+RgOpMJ0dBHzsYOfVBDgvNvs02+WqgH1Qkn1ZKlHMQKDnXrL2
ZBx2lLsCm0vxykpcbO9I3RLmw/wHfo3YPBodA93FBxzs54Q23ZCYGyN+BlOy23AY7eVWCGcOyZgF
dWLtF1hSYsU4ofp0LwiZYprnsLnvtGrU07ltTpgxJqp0rk27Loiy/qr7oi2aXWggBIDX6CkeZ+n1
qjp/BRBDe1xF0+YtQB4Qf7rMErxW2aXDhMMAwu8E5CHA4uiCenM0fz2l0TG0TGHtKWD6YyNDbgvv
SRXhjU/o1Ur90Rs89sHblU9WD/g1DxpvOVIoSuIdEKmFRw1Zm1h36TiHjiDlo7XVvgkrkzSg0oCh
fF/qa5+/kPeNsZC370sy02xF1XR7CgqYtCVWmT/Y6UGyWUuZZICV5PD2iTpOlcBoVKhq1ynmwdOM
9pVOFd3ZB+1Rtqj/wgtHwO5S654Zan5278i0cNT8QL+nvFOPw30TJ0dHiGyubKwNFjlUoa58INjt
sjjN1oTu/AoACImn7VET4osysMlH2LrvYAxBbuHaVNZ6gWdi2JKILeOlKVhfm8AOFUmfeC2IM8G4
Xu0bGyops0dJVUttmaS2AnMnYlT9vFiybg/cWTL/oKsfHRFVzbLAt1xTiP0fsScOcgbZ+9GE9d2i
91PK4eS2Opxkd9vioPE2qapOZa54RWUGdYOFi1NhyaxXCdrN8vkeL+VuJNxle45pNlsQTv4ksnK/
ZEVszIPC6tLR1Qbm1d3qUT7w+0Ml2ize7NpBwp49GJtR4QVO09cEoRCVOEBr78fLOmQwzRT+e2M7
yXXjkhIZdctgCN8rH2P1dKX9+uja1MUxswNoWWDbM2AMdnOF6p62QZ0f1zcAwxWSNo8nFZzpYDq9
8goh6881b0+glVCUqc0Y3cftO0hNgI+eP0kmley0MK6XrcaJbE8va/ZERvVroPD1dHYWZ5R25Itk
jupxxq6G2vC5Y/wSPnro6oR6XvgIaUqi4GGDF7Y7XIaVhtlSr3B4LUOa+iVPLO48ui56bFM2n0sN
3gBqZE5MD3c5huFmPU72H9uwJAiuaNxYoAovNL+cXSWbCRiuh26KRRBFiM6ZGTcPsuqOXt3nDT/I
WTWxZLlpzsmCr3dd3gcBFqFSbvf218Y9wKdHY+xW7nU0u6Q70CjPQzDA2ZN5cfp50cvHK/AeRvT2
G19UUJtMfdWdYocem9cBouOFtsxy9vDWzR7E8PhTWx+raEF3hO2iNzhEn9OMrYhYyYjYMhvkI+H4
lVm1BU1X+c5YW8Ek8ytyvo0RwafrUXPWJCRfdmIyWUZxcjOVkG6J+smHduXQBG7v2s3BVgdAEyvt
eYoLo4M2UUBNm3ZQM0bOi1FVgkU0cAzfIyUx7Dl4OvrF33NISUYc2gVQwIJey6hIDgkFNe8ti0Qh
TYdy6rphxeRTCQMrpGjbelLNcU0V++lGuymQAuVuzA8oergKMBD7tmcYHJF+19f7zsV39wYX+eF7
cPkL9BLPMiDhe3QNOvGx7nzdvEYNatdM9OQ4loWfN4J6n/M1PHET+L8QIgtIlJrdp8MBE+7RGZyF
CqJ8PybgqVPlI2ZfvE6lqrmYdWOM9qdgU3iajwTHP3L48ZpD/Yp8UwIq6Nx5au9FeF626OVMVfgE
vfcqxeuA9Pbh47zPfTNSDxyL0FsAxuDus8gj13Ak2i2S4Qs+gLzh3FmFgpmglyK4nby/1cVQj6JD
5xtjVqkzGW0PY8ij3IquENnIMtjsDp0bHe47/PsOXZQRoaxzrdGd9lkZPN08756f1K1YRjXqE3rC
Z8AOoi5EUEUPhp03shBV7ExHqj+OMg+BU6ptqG0D6ksbeUK3MUVR6ATK3qSblACI0TD0FX4su+oq
ftqrh/aA1KlYx4SRZ/mL5msFLQtkUoAEckb4+TbETCqCQRpStS04p+Lx9IGoHwH1xa+THtBgTH58
u/+X2mf36l2Y2MqK9qWueBf5dn0YWeTHF48Ht09tbk/U6U/9j4fl6rUhkdUDjRPYbPzganUQr256
oiM7FtkJ9aoHDx4T8SFeDynrPZf7kek9PkrWH+nUtw9i2fdW39nuFTPYhYnLPQHW3vtpZDG4ZSCA
GD4uSDbzKscvIcu0DxvEKJheHu89fiFl/L9wUJGSNfvLlQ06yXR9dQ917Iw9Hi4FI8H+fp4v2aPD
oCV0ZxZJEQL+E+cbTjjmemQRm2gyx5DfGqUI2VZh75cVK6QdY0E4aaoAqT017GvIodi0pyrdug5o
NrCvPePsFkkEfGwHgRXC/DxsMWoacDAOjo7XcEHxdh54TA6H0bKPkd53Y68G0KDdOZa9oL7wFiO/
7tnQFxqTUNU2Rbm8VZSqlPJndPk/jpzLtxhyTA4KCOztMJgnbyyvkoUlz2ZI7hA40OI8FMBAD7nL
V3qLaPdCCR7DYUma4pImgrO+0RlUhjHO5UETj+0a6kpPhztw6qvHCTg7hIna9ZB/ZnjZxanHzbpg
0uQtsTD5QrpaFKdIPZkew2jXkPPDnGJhM5URxdWnUb9vyDlxmTaM5CtWvaohtKlsV32AHKOavZz+
nBFht7eUFDeoa2B/dhRoEoGP5MH+5DnkqzYu7EgES5E1JctAY4J8K4sNCsgNuN8O5Pm40woAQ1oe
IunYm12o1Q73MpokpurMPIGdHhu/cik1I09Ch9ul9ntcSMKd2uXX5ExiL2fuHinGGU29iGZmKTNa
uaj3SmHdGhw/T0W4ZEuYeALNV9DxSz6/cnD0i5fmKGkkUEiLJjJVo5ybb3KxJN/rySISrl9ojaQi
DxPqcfuO05djw/t+qcQygdrWqZWFitgpT0Pp104x49554UHGeQfz3MknP/LzPGCpiVrLN1nFcYr9
N7uOr54gdscupn2wRGQV1wdLgDMvWsAb+iG7iSP8BA594qJwwa5sSsBXD0izZzF/fMj8ea43LtQ4
5iGCLmguTsnclodsUPhpa7JX8DhiKVJHzLHZN7qLdYvoBZPQdl9ZLkTvks1h+24X+U62HEkE7HtW
8B6ssNbzng/HB0u8LtznO28+JzjRhMjg4JC0VU4ftyt1v/nGxe9+tm2gzjWKeiGk0Zv31G+zi0AI
VUjIAMVz8x7/M3HkPrFJGfCeqWWe0nFeGgVT8gJYFLfV4VAALqsfHQQPJ/dQy1dqAWgbEJXsJOp0
QVCwQOoImDxCrjI0GPlif/HPbcDBk1+/xNatBqTVMyQsHKlCyF4wTl2fSd6YrfY//JmQzZRB4wxD
Ku7I0Eu4Bo6JdZLXCaIhHwCog6L27tpYb41sg0br9RjW77uS2+4FK4MbLprvRu2PkcT/8hlcPKEu
/XYoRR6FJgX6OdTnjr4TGGFcz9+OIWqApGQmIczqdgdSOgGTnwRv5pRRaXjNfVkOKua4FpniNjwl
HCavPBZk3YHpWQYXZkEptgJDngCEmwK3rgjHwdkKefLp2rRnyuJxqX934/KouNUkFdulBRKp34Vz
CuQRAMBr1UbpsoK5Da3eNVnTvvIBduMXjukLMZ+YDjLt93kr4DWjlDU2L/GnulqNShXw6p/eLj53
GoJn3mh/w1j56F9xbLeDzYTIlsI1Qey0uEnyqo6N1bxoAsJKqYl+lU87Cbl7PSmaz+9rNphgvuHN
Ty2SbvCSsp4M/tGb+0Px5fImiVLr7IA2CUgp+HAjx8uYUFObduhA+YVt0mJe07mqy8D8jbcK6SJA
5gCDue0Sh4f5AjirT8fC3fhvx1WzdCD2F4n8xs7J8Xhy1pOui8BX35bHyiQsXbdNbRwAUF5U9TmL
qB8YvWdNlUQ+HT4U7Z4B6V+Wj8kRi782Hg1/0CttLGIHdiqxUgs0xlGz4jJPxUZ4/hEtY2VFT4eJ
v1YEgFXspmsefl6SjO/VPdQeaPh39iNaKwcrZPTREDeXKdHHrR5Ouqk1xM3QdX9YsxFcgqJsrZUc
1yC6TFqm3xwssFMa3hKnUx4BFuD2iUq6l/fFtWFMblo0oMIrm3320dEEPN6d+z2CMF7laF/odlDx
yjVJEapHuvOV//nmvjVVl4KoClLTJxG/y39Tidl0LlYTXbl+jqbKnvBivHnabUkofGhHR6kOgV9q
EskuW+Ruu9Po1b/9F1aXkoOrWLDDIsn0PuHAcfs8895VSI4BK9pjnYdv9S6TawcZjnyZBkkXAv84
j67bS1J23ywraWONA+ixPfjBXi77liw0amc2akP0jwQP+4VCrUdwvk3U0Ii/CXXM5DVoghJ59PjK
O83vEAnRTlwfEdUKxUTcVCBFiW5xzaMCGWVO2FSXkCjpMm8jzI6DAiiPLw6oNiKgvoQisykXbTT5
TnuG5lUubyppKePQYqGK9L+0qaPBUf5ClbdcP10vnBSJRRY3LTIR8yqYZfGk8iuaaPgEsqmM6XZP
PM1MYLe2uuonhkaL+QEBdDtsKLw8pZghzMYEzcZ+5KwaxmMEhaHdf2PrGFoyShw0q837MhITMHme
iOsD7U/oLqfRFuH4lHZlCyJlHHGb2Ay96pVlGPlOMikKHOMFBoCINyPQ+YtsR0iKUoqFO9wobd4T
/YWcwrqrU+6e+R4Xpi8Xja2CF6kANzpPwRuTOlB4mIR4SLldcLn7x7Kc0PMfwqplWJtkXdLTwQpf
LNlw0VhQCxpLfhvloTGHG5bllYaK4dgY0XgoARAGbXnK9bQJMkJCwCOv/IlzzZFTdklDclnCI0mt
faIDUyksHFjXvvGmt5n+sqpSGfdC/7tfm2wzuIuA52FkmwyGSh5tsDEvzq+7tf/XSBSW26GeMj/K
dldiswud3PAwBx9RFdnYh6qxS1Scl8xnyqHlubTPoSrJvvhlYWM1nFUAXMvurIs32bpEC7k6cegL
JN0qF9hTqgbGg3poCny1oLwhVjMhb/n0yhaWRFjVEdrdGN48vVMV8IfiDZF+PkXVA/ljEIVuMKEA
jdPwqTkvGz2J1tVzNBljlDgKM8N/yWUKUNlIR25BWEOcNR3bcNO8erX+WK0lMQ+UY3X6mJdjckaO
3zGtMw5z7bYcVPJY18OuIVr2lQMD6xrqqb8ljPPfp+Pe02XGp3NHl5iFB2fisyJ8deC5SKehSXDd
kwMz+Hr1c5kcp8v6ZoVLjG1fae6bpSPB3BKpNSmccB76tJ/AsKv8bTlawsV4gphhm3RZyrXABGua
kwdDmeZCAQcsl5nf+EUQEALb9x7QjheS7xdDjaGKVas0r/IpV8uhNnvw3bfBgYH9IjuMdMm3LCTE
YUlDY4t5D748j4i0iMmSOx2Vtz0kAQHd0sNnmIDEpqlvZkdmsUiKu9wCHEGHHghcsl4fjT5mVOor
vTjfVWmfQ5TOUCL8c7hCJQCCXBnxNOBRd6PSXvK2dlEYWmj1NBQ+DSTbdmzgHUqvGkKsmUe7NI5H
HO+KNdahZ8y0peQ4tDDpYXuFLJLxpiYRadB9cM55V/fur9vPczdXTuNd2eVEgobClrVDDMmIQ/g8
5P7lW5i1p+9ea2nCG+u4Xd0+D0/NKwOHztWPvbxyQyEKdPeWmuiXCKYGK2cOG39yj+4VFLkqUWLr
17TNs/5lw4CKAI5P38uQVMFM0NmzqnLoFOqg/v3h9FWxL6Ht6kBoMPth0AxoXySQq3HFP9QDPNJS
DKT/fXvlzUkUWtHMxWkhhq8yVub9fBzwbVxi0pv3cw6Fl3myvFnMFD176VQyJ76HV8DdIXyBg0+V
HeBE6f4IId7qIFm7CE2hvCT9exP1Mkp/QjmpfPNLXk21ZuTbEQtaFl9MShha8onYjwKxVquQuU7a
cGzdThICcdOa6OZ3I2kT5UcQuDSCNktnznDL9u6+rerW9gqtzRMKJZ37cUEQUDDjva6dJLTos8BW
3SHZ0I+VKWgbCWJDbJpW7dUVJ+y2KwLt1SXdMOtfw2VJPAQPswZN3XPpE7ECwE/muECUcz475fO5
c8rbm4t00D+idwBymM4VO7hrXKsQ1i7YTm6cX93yjQXuDWubnrT8W2wD2Hu2WmFir/uWBQFr9dHE
B4nVII8Wxp2/0Up9pb/4Cm3jBnNx1BaIXqxLzhf1UYnRrljd35LbyBbsBIuG7mT4ncgkoogXvxrP
zZxxv9J2y2ALuXZuD+vWYvYpqCYATXb0dFFtxfmmxHJ0XEpAdCkZ82WZP8xfL5OY37tUt812wUnZ
eT4MYTzl9ZS9AW4cMZXkyR6KF1Q/26VerVWlVDhjwyWV4LBD2VAZw1/6zTyxtCHOkodVfTYxhRhn
rRaalbkucWU4cqgG5AOCnEPbFP8AwyQbQ0sC+pXVKjHrD+VnxGXDzcUBJuMOpT9o+jEX93EArdP9
RJ2clsF0MeJkMTpurHFwJ86ru/1dmiXZ1yaD+H1GAbfaBfRZc2quw8oWDrv0cQZCrEx8KKpR9Ptk
49519w1UdlOaHWrqzk3eCUD5wwXXD0uYr/39YP5X4cOxN1SEmLYFd/NcUJfmj3lHCFwcumOgPLBO
zUTghzZbQDW2+stRow2ZiuiD4pQSadvHq0mkvfkqBD8AzNMoU51QWEJVhHcn7Hrf9FPgUNcErm9T
mMvy0GfwYiVxYwSH+0loWmeTl7j6l10ewmcY5vqkEO0brewSianhIw1on2gLN8g7WGmQi1cgFakk
tV94PlNfGuz1TcQT6fg5TIUQHQWv12rjukuFCwfkIpNG7Yh0kPmciFMk2T1Iysv/sLKgxpqxBzWK
spm78uEEzds3SYvPKgMEza7vOfHqqi0e5ntaRxV6t5FKCa+Ajk9y2+DjIvRLso/z43yfFG7BJ1za
RlRDAYjUtv9U+opZ1R0ThGNMhWJrmY1OvtOClbe65a1ruN/tgR9i9WisW1XBz6FzkBg5jBvmzRj8
2l6QiNwAuE/2TaNoSUpMrTbQrfzudG5O5XjQ2AqzvAMElqPIHIJRhdwsG+QuUZ30ytcuJdlBmLAf
bRwnPjC5XEvCyqrNW/wl9osXWAwLzRLHQnZn5QTqvOyWZQg0S+8jSZH4WSVJc0PzEz3AC+2/TLln
wnBj31yY8NmIn1IjiU8CGyWW4PdHaK+WjNQL7J0k9E4rMCVq8/9FPtt5rACCpGF1pEHUy9fNJ1RI
a9uxKEjUFRTBhRKWbt1fixnkKCo0DIIh6rV5dqAG3PrvSu/LA19LEO1PBQxjr3XfkyTMY/IWpo2i
2OmewOhcIiw9v/+ikzqyvyf74QzFMvsTyPjw8hplwmsk1oNzal/a3/c2YiZW7AI4oEokv89wKFa8
c+1ortcUfpO68Wam/oJjcz+0JpUTF+Lrj3AFJc2o0IYQxYyI2ZbFERFI9t+ACo1rt7zOI8TudMhO
WDUNsGO5rF3Lz/sFHDRolwpqTJwWPilBaGpSrjWxLYaDaYO9Lj0QpFhOMm8Np1oSjB8dW1ASXsdG
TRiS2tht1nZ/U36eBCGdPSSqk8wRG5aRZbQo7LFnH25GP1jwwFl98WA/f6Qe6sFt6T64cxwXSnJ/
RMqWYb6nESdMvr6YR3eABMURdz88WJ59EXNLubCEkV7d+plgAbWJf5J6plc3UpItqxEsqqjdh+76
sT7q14QsqBsinof76IaXQ4VP44fzWLuGQY0+driQYYFVMT+Vl+9MvccAYRnVEt+3HCW4cobDoDAz
knXmzNhr5ovrMTFF/AqQTNrwzIO/rBAc+Rphag2C8npGCPL8FFsKHoH/V1zWnrAmsFgSpCKafloQ
7HBDD5HD9ZN8v7c149L0S1LndkOxGkgtzOr3verzR5VDIye0XAjeaLEOvyAQbFw+OZAO6Gza7dH9
5f70si+KiAMb1FyYsesF44kfpxxuMspTFfKzM9dLnbM46i1d4O8fuMCvos38P8sqLqAE1lefGHa5
q2j/zgdpt37gfDedmon7Mm6e2NFT155jO7bNBaxvB4b7mXhlRrShK3jt7yathPBQ6Y5+D1oeEiRE
Hf4vsMnmv95mqvJJMKEvHrvQMYZotpapwG8VcIuKWdyw4Fg0nwLcWw2h7nYmc9b043nCs39U5JPo
9qBd6w195P2jV/f3RMHwIaR/JQqejj1jp5g0GMZOmm12HImq4NZISEbX1zvpYruLOwQDmIwnEEIY
+dLXGrCRXjpKVcF6p/mLuMSx3sjYHVP7mjdrWfciuwOHOOjQ1w+kVlxMLfeFT3m0AM7PPaOf2ZPk
bnMH3o4H7cpSkEJHisoXHRvsnY5XxsaE5YXSfPCWL5jR+N7VPYLHWZWECNRg8BMQyv4y1cWFhkju
tinhSR+fP7DmO7MAhfYcEK8GM/fJEyO73zMri3wicQvAWh7jZr/4qByh6VitTKAqEmLEHG8WqQ+O
OMn+iX4vqIyWT4+3zIUMiqiK7lQxrKNjvIuUgUo+IIPdWQEI9IxT8VmZMAM55kM8grAETorIJ8no
PGUUeyh0LWcbYfpZMKWh9X2/d5djF44JHN9CzkL8CE0LtXc+0odVAgyOlglE4OeyCE53Hy7Z589J
KqGrxE4IV7KVSu+tL+HWWSv0dkLDW5wUv3qqsAtmToVDB3rUSvXcU67jbJ+ZQ+jtQM2ce5xXtbOD
NhxfgC3waJq0LP9FpOsIiAx/Tt3Nda5t5KWvKqbtG3zTIthHS4GJaSrZUz4rYWej0oTOZ/T99Xnb
jY6BAicGxbm9wGUQqMwyVttpqJfxjd//C982I6ufRIbDIaDexj2HY/W0P9ubH7i/ccjfy0E0JZ4F
XELZQ/v/AWCqBFBtMYBllX/mFOFhhQKrbhtGhI/KRXGz++LrAyfgbhHUKoBDsgLyq+u2wsKkUchk
mB3yAQ/FWkQPfI1GoRu2mYQ6Dt2V/uO8higQahhSiy4KPK2G6b4BtYtQyDzElMwnSdg4I7OLZaS/
LHrgi+34jNn81Y3CktJnj2PR6wMkzmTWu7x1GGSPhu7PvLAsPB0Gyjaogr0dPeDa/iZOEpMaO0ms
y9nuOxQdpVwWlHdIY8oDE3mipnkyEqSPB+2XeztenqDZ/5p7jtP643o7xeOZtmc0cC4XSAsaJXab
Uw2/nySktsiHTBVB9k3IzdAx72mC7UOOuwZWenlKxOdaLlOBD77XkIjE4msjp0XRCzLPirmDL4tA
B1pM28FSFmwGZOKoQpuhP4sRB2F3L7c/prAZt74euhaGS+9KwP+ACmWq8+I8PCu1aS/SwO5fTSfU
580/Z4F/7BHzB64HVSsUkJZsqsVUj6hei+MysgC2+EECcKvypbl8ID1+ethBbVMFtlM3pM5SjfLz
SGI4upvZpBWAsgRfm1Zkw6U0lQIvv+KIlnC07nNF10jb7bKLNJ4Aicet81P9nxu5di5RBdNJHvyh
NiaiL5EizOMdi26cMhMM/+9XqAF5oz4wsPAef7YWCAXeUdIXjMucJ9bfLwTrBEkPVH6DbbBOSfD0
/uwcKDdO4KBk9N3mN/f9QSbS8CqQTZTrnBALwr2682YtTa4EmqEEbZHApPILqABklhY3aGdvxCXL
tMbNiZ9SswuS7fa3VIIqYRbObeE1Q1h2Y6XgVg5olfNTIXwOwUbAS+E34tyUpiVwKjhdEXbjmrWk
sxSOHPjUGukcem4b9AKfQpYNcvh6HQxPS4RSGxGKttk3v37nwRBq/1IYDT+esxgmwQe8pSfOBg/5
n/xuX20B325zMCK+aZGFobBppQdgK/uuqdq6ZL50fNQg8Ck+ReEVxqUkQdSySZNEZRdddH+TwOBb
FPkJehkQaluwB0gePg7ILkjV8OPnhzFpmz7GUMlZbzxVrHV8PVfkljlgwHGWelab563mXVpRcDCk
UuXRcHxvzXsoHZWIroV+KGv1zCqkqLA3zmi3OuTj+eeDhHuoxoGtqKe/oAs7b1qMoZoWtYY8/A2N
GbsnOGdan8VseFLZ+wfVlGGMzwL3dNH/bxsItr3F5w/pVT/vMEGy76/Py3Yi2bhQdfApcQIb2hVD
tbbHQe/siCl3EO8bEq/aazlhSi8hSl996tHa2bR6nibuO6pRkjxNHFku5dtp7x6X3GtT3kMCzGpP
zPxp0xe5YmdnvKqsdlJhdsqGJtMFeYNmp1B8w/ZT5KlyNLqSbFk5SGprei4pXUVeRTQK+k3074uL
2l/5/OwZWOUpswy5V+HXfwntWOV6eKIXl9i2WWivvKrQPB6SK9Hsd1I//j9/8d1Kpq7Fq3KWZto8
1Aoa7RGm/22EoNH/oMA/DSF82RVcAzUrswuvPEzr/3iFQ1ZkO6LLbYEAKJGDtWbxwfsubIxMaWAs
VEgUC6wYx3WbglJPeST1PpdDnzq5xHW7Adhk0dj4Rz8E30AqkP9ykQgiyISzdTwGp6bnqapO0PWy
uETMhG81QZoj1S7NBg5eP6f2ja2hGBSnMpAVfvBRktZSZpVVnVxrBEs71S5Czr2wRcRKJ0ay8oz3
W3voMDJHoJDzcJTz8JmiUItjknvE732TdXT16nJK+EY9uZXLdz4o7lRM+IyyuPSGQwo0A1YttPRk
9i+zumxM5llurmp+6A1RuFarxT9f1NjXysHnKb/jILbsJdqQrJH7wZ4EFOwOL6TXV0HxIx9nS9ag
tRGT4I4FHJJMiExArAOO+zZwPK5vrhzZmj+2yk+o53qcPLXmV6ph4xT6kMrWHlby+ok0HX8wVXBe
CRP40abanz44m70jAR4AISSrXGGehNkUMugS7L5UuNJHGagaANGzPqRJK5lDNnUMs9Zgywor/siF
L9v12y/d0xJdDibH/WyKzWOYqzo8wO0vM4HSKPfIbsPOgEa0vQqTuF3TzLdYeLPuMxFPQv2DadXN
4R4p/OXTzLhZpc7GnTENa67q99fsiuOYLjEYFz9Ux/Y6sQ9bw44UigSSRbgQAhnluqqqc6EPB3X6
evVY3cROVBFkN5YjM6RpyzxqsUurj6JL2OzquZ+AdkiWXnHn4yw8VpuTpuELaVFIjQw0f+/bZcmW
TxgYexgfqnDJ78MJLQ3lyGOHu/K4mbpGIpJaPaorQyTPpffKe/8oIBmEvsuXeYO68wcZAiMvka9W
jDJtsGlfS3T4Ix7/MxYs5wQ7bPZ8X80ZkKLyyToPnHAfY/Mf2J+n9yPflonOGsdvp2tiWCCEjp3N
55KGXO+5MYCsZfwKrBm3DobAVHwuuy7dC+IL+ZXllVV6YPqRPKggq/eIPrgIjSyEzY5jCGjLQVrv
CiFoStKevbHsKhzGUeHYBotCPkkzkE6G2lV+qlsUMhqIR/A3Gixvj0qn5ooVrwHOpHoaCFhNx8WM
AMTFlm08x/GwUt/trtcqNM1d2a4GNfEGpCWiB7tDHSt8CA46xBbQUifae5UJM8tw+su+Lxbwybd0
SQihnhf63uzK3XtYBS+dRJUWarhTG/Tty3vgBo1A4GJYhUGCcpAqNCsVkDQPxbgJUzAwMXhsnOFS
R8lpYmQSDIsZC2z+GqBlA4Rcq8l7dStHONafRLFh6Bgl7Vtyi9upZwzlqvKI4dUo/LdLqOLloJ+C
z0qPLAHYwt8l7sKNyLhLcFe6b6RjuQzrEGKrtf/z4rUJGhm2b41W/Cn1xKLGMi1r8Uhbd9kYqVMY
BIQ6C7C7Q+Cgonh1UKm18edWKo1PASFsdXEVAs8FCnOBj3sPICNMkiTjlMmdK0Y13V8DoU+l34Bf
kKoNHTYQUeUdkK5KfZyyrJYdWjMLV30nU0eCHFB7RHqJo9OQm64q7cHIGNriFrCnE0i0zSFSTaWm
FuPG8kMvMEvLxVwI1pGV5TCeF1bwFfBsRSxAFyNTQQUjPmmzOdn/vijqvjfzvwQSH1Q4TKPSONwL
bU8d3fOobIvg8/7Sb5+0ghMzmU8zVxqSxU1QEKjlF2zwr01IQZFQZSSemCXaqhue/gsH5JGOiqQg
bbY4wxrceIUC9/No/IHuqywJMqKWpB42CnZ0YdgNvUXzVQ8RyG11ZoXYNaaA23W8xCYH/ucp/VW6
eJxYqd9rDyoN+HlX5BPXBmV+ADuthZSMD3J86TMAWGQJda//3Lu15JSEF6KOorK9BIjVNBTE1PB1
EJg7dTQlwV54DxdIfaGbptUoCts2bIAbWwcyFZ0viTz81/0TRbY3IqYslVlkuvJF97ytjpJua/wW
mlRsMAhbZoMbzZPY+pByOAoh61PysAd8Qr1z7KXvR9FcqHR8i/UQLlUShYNWPJVKOXb3hJNv8Gm7
ggGSQKzAOLb7KWiE659kqSvKqMPOPr5ld/dM1gg2glpG4JrDuoQL2ugvZmwm4P/f5K8GQIkEF7Um
wmF5Lb4PSK0FSPkc+AzjF2hvK/2lEm622RKCAeU2mz/LmpuoqEOimSoGZ/VuR5e+kzzis+xhpMZx
PfV1r8pVYwvAvixPKhhjKBCfuTKqgXN+tG/vkBAdHoOEWhNUzZz56pa3mNQMMbZEzwu+uz/N4HS9
O18RU2LI7IPVL0Hc6oZekVsfNqSNNZ0B8Af4Oa61Cg1Bn1EK0nhXgo5IHCDO2byaFyZLlgXMfZoX
0QdTFYP5EA9ynlqnJGhdE+BfCE+NDe0pPMSUdVi9J16TjLLY0ZoeH7Ncreq2QoY2TP7DZZeVAjSu
r+vjOG+NQYLenfMe4kEjNfz5UcMaRygAsOZXtZAt1Nsvzq9/nS9FtkS5ZkhEJoNDKK2178i3LlDw
CaarR3X1pChmoSZDqXisexzIhboU4SiSB/V28Us+v6ElqlaNIDgRXNOsHfdCpI0P62WOUHa+wvqb
23ki/NyeO2l4nhiFROaZfpxeEVPL+GtOBHshz1nSI/4w17dNp16FVdEyaLaV3LPc9Gft8voU/obl
Jywt76JqSH+bZwdYjQYHKz32cXd/tAeFwI0xcAaCdNpGitPP/2dbEDeBicjGm2dgJBUwPbBRiH39
gLYsJr/XPSKD1arc7xwcxoYqLjCl1u0p0d7fdqgQ01BzvsKH8o1d6JWEkd3GCLE+8IjJkU2z+0zb
Qt/Xmp1rp+WFNEDneWbYJMuZEc+XZrgp69BQp/WmkWNWZEv4djTGixGeTFov723sY33ibaLAm+X5
lhQ59Fk4cG/s5FHP57vEJFnkVHSaSxarSy8++rn65iEIH9dKWnSJ6P/eeiqfeaUz3wDrUOKMIFHp
wC+48sWrMPYKX3CfsEMDKFw8tyi+KZ0CQE2Culhdiv3H0UlWn2sZXkS9GKdlFqVPZA50G625m2dY
1SaTTSqHzrvc4cw7ingdfm71qP2HcFwfDLf57c2WEi/2A9+7SxQ7XtzUQ1jQHTAsRGW5pMzaSXOb
IlxnXedr5QlwOXpd1+q/2sdky5SQXZZgj8GbTkZbq+MtdkIDKF68wJzrlD5P6LMmOt5kIiSjSKn1
Wf0+Ij5YVcu7U07WTgCh12slIhkvBgtwlsLHhMi9DxVp0BFjRFBSAaq+bBSNbTjpfoHgHAZA9aLv
BF6XvXQ9wGJYwnbYpYTeExHXMD5yWMdzFLetucyFO7stia7u8SUj/fsTJo1CeZ+ruhcVEIW1O5iD
Cx45APySC0dP023jQYIcPG+eHeM2jRdjVNYfzIdRodqXvP45E0WgCwI6rdE9EVN9PHJx+lDk9Ul4
FnhivOY37VUeKQFoGvOJT7fLcsD3fq0vfscHw2eIYbKkJb2uBNIf5Hwro2MPknxOhTMwrOxB24kn
AB2avKdfU8bdITmdB6A9XSPk/HVD+qO06D/9wE7ODbq+eAowhAIWwDZ7TZyD+2Q5hjEi5L3QFwhR
AaY9FNjUMcCScClk0I/jCyu1qCQxEuGJR1G+M0J4uoHHdC2Z+o4kdVHLOanT9A7zGi2IlvajC5u2
wnb8kxgqbVMfwfa0anAzz8gctVk9HLhGuBN7y9rpTRLyG2cKRlyHO8GvGX7DisLVbXBQvwPqVB8j
8uBu4b5rq53S3gVxp/LZjEImo334EB9OXK+NL1qNxeBsQKHJcESnsV1FjUg6jCQBn3R5fNMmtYct
wfHdkvZmlnkKB3UPwFikRSkrEgWdMzI3iaNGTi1Pilg6C3QUEYxNH81uwc3BAW3DNEpQpYO1J5wz
LBefp1Rcp3NqDu6ubu3r2E6XeGL4WRbfsHNB0T7X2x6kIiJfAfh1soywGuDXVULiEz7ABUCYRO2z
LodLybPLT/otOF+jQMC3CS1b8wn4rdQcOMNq/F2x/1hla7CrU6PGVMdyP8wVOpS7O0P2j4I7AGAj
8GRSYKJ24VbIkCSEAXbWga2B6XxOQRbwpIVjSXr1FRmY5h5nU3PFGmnKgGrioyYy+pY83fIzd/Jw
fzwVslEA/pCw6O++FvEg7hYXInQlkCzSOEqyrRBi0lMm9f7ZAYtsMf2rfRRt2HOMtGs8GceuvTEO
hv/hNphocJeATsZVQwlEC5a24ituQv3aeSFL7jMwPQXdtv4a2s7oeUerPTN6sE6EKIuxueDKOR5r
1xe3XIBMJUuy0y74k896EG9fVuUGa7hzsjxedDK/cxBr6WwhXujHOcRf+GhFGuRUVoGdA/sohHto
CMIcb0847N1ht4GSn0i3Ci8yRLBlJ4gzaMm6EmgX7YWnsRMVX9LMKZyUq91w5BYJ+KnWNw3ZfnXw
32Q0tv7u1DQWHyYa0RRkdHjFIPadgQd+yzre7c+l8bk31stp4yAApdwEP70Uwadud3LbwvJxCp/P
gjvflTm1eaXPJZ8bK0gat75kwOa6MnGw92Q1iL5ZRfyGJuq3MkvzrkwfzPvsC5s9ZLIG+mipx9Lx
WKKy+JqW+1E7Nq7ush7NlsNDrSxgUr2w8tObl2gpeNFsJhFuffroflbLER2mIO0wSiYxv/y7ujMb
ZoIMjZrTNqEO5IBx8Uu4HQr8SSS8KmRANFUKN5bR0cAX13gMukfKrkQwb0a+b3JzqUEAviAYr7TY
ufxDVqLFC9bMRfu/Emueu9MANaa/TwACB08OoRNxkxIpKj0DMvuzh36rXx4ttm7dqeO1WJm9EOfD
YDbb3L2kkkLB3l3YK/BEztZMtOpFqqHEER/K5ljA7rSUHKt+EtfFAQvgQL8qyb9dWxmpj8h8U70+
Es5DxpR1JWKkn5NGzMnzecP+aqR7k+KqBe4sowfFfNhIu4UqLaF2cibQ6GBCc8/BoxHdJcskqv+m
mMGQhY2SNGe/9oQHqC0iAJPXdjS4CmraTMXVRgrppwXm955+n2K/oLq0TK7+jXFkvJnfPWyAcBVp
ozWHpwvraxcYAVPHLoOn60HN5D3I8ev9c0W6iVKPIKrBrJpo2L5/cusiLlJipKIrXO83N2QrpMLx
0Hw8ZuSM1/EKPt+LZr/91xXfq/o1k9kSS9vQ2X0bk+uc07Pl//eJYNVL9hcBF8qjPPDCTFh6U+mf
E18W+p33QIvk68NI+eubHrKl4/aElFiiSTUQJTMQN1nJvNfT+6iKu3Clu3+wSDfjtXfL4W2OQdxA
aaxPOLVxYRWLWBkyolNexs5yxex7kyHksT+ISvE6lbMGIOG5xWZDPwrtSY15bKqZewVKTOkcH/aY
vf0hiwNtAHlo1YIeW15AaLPs3qG6OY9XqtB1wvUnLy1tOcf8YC5SHA92auj0/btumMSc/PpZULbG
0EZB+CM4hsaYWa73pCHG9KPU/MjTlLBb0Zfp2y4tLGZwS1MuS5yVpUyKTXGo1mXGC0Rkr+rCS9yj
3NwNi2aNKGq+u6PHaLCqVewQAJ56y83TuhldFE6Y+pQ/wy//J4DZf/7N10eHxjD6HLCd8L+4mR5J
CYjI4kkmWyaw4OYZV6vWhSmLV4a0HBmHrrQ7tTDlv4jCbfCjDZ8egMiDVwWLTQRezK3kRCQvh5ix
+39ZgbP5R9x/plRkHXDmHv587tOsDiNq/R6fsAqfQwV/D+0NEOBm/Uqrq/eAy1sji4r0Un2lZcDQ
Cn5ZoEq1BmcRptvQDA12eJS/BobCUIAK1+Nm/ZmTM79988wN+FdjEb+H1FxEGHC0Vs0swsr07cft
Qnqua9s80zJd4TGYfhngvwVnA5Td0M2xHquNy9xpq+oTkKv/C1HycGQHN5mNLCfhLqC/HOlXIilV
DqyTmjEpUD5OqWo/ZppuOhXOWRTafBBZ6OcIgz4hwKfZvMbLamn0aeE31LydQl9dzXvXteIVKgkQ
s5zH/NkQf0KevPIyMUoQ58Uq2kJaQzcr8F8LIdE1ActgVPR61KzreOGEQKCMiSz78ezSoMifaUc3
OmeoodukdKzt8TI+RMTdGifWYe14vUFQkOAFEeiziGWIBtmeql6ZeUy5QrtIX7r0OSafd1OE9b06
eFO3jXu+ltwa2uq5iMDeSyMKizNtfjRxMM8v+gz1WgQN8N5tLfV0h+9eckp2QOGoFOo5skHLzrU2
UtZngHvQ/0UoRAYbD241YF5lTeBodc9zt0tjCoVN4bccFK7MZeTqCPrmiUrxbXLex6DGWlz/SHqh
hGTkNzjOrHDcWxgHWF1EuT3HTkRzgJNOjgUV8vnpPbpx2DdOcooEEAGt6IJ8jF/DszrrCrMqevjy
i+pfCqCppg1yzjCHiIheAEud+Q8YfDiQcd6v04mjYDHDHvz/RaQBh7BZZtZvVPLmA4289H1bt3zc
XlGwtDIq5SdFjCQwmURF7BMSUD8uZUZV7acCz37wF2bRxZTLcR1ABv0VaykdsfLZIL88TTNXMt1Q
1nBuSDk51Fgnu2IRtTFVMc0eLHK9G7duNiTMbBcO2Jw2UIJQbfacp5Mi0mmklUFAHx3uPq6uEbAQ
O0U8bSpffs4F/B3GxZi+DnpcTyhFUnZnUGcGsCdD7CEHQByXHb1ANhBgU5y1LwJBFoIQwBtXaAom
+IyzoVbwYDY1yBUaAAcxH5gY/M3rZdQF5Wo8Wb5CefpOLOC+ecwBypFHYD8oBmKy5d412u0IgaA4
/IJbfug5Uzsdy82hHQ2e5ijIGpJXUbCZf5mnp0pN7ylTx+EMiorCSQ8iEurjAw4FHNgChdiP4O2v
o8Ujo0LvFmLV7JADPYZA+ffiUrD5AcVgQ8Zm22kujit5yWgn6oTz2liFQ59ini0zLyaksebxB3Lq
nBpz9mfpiR7hTgx8hgnbeeuBNlh6YGvvsYpH+e/atGpgB62xRU4bj9L39QU4d5tUiQbfMcf8n7mA
qf/bjdsm2TTJBv9HdugHFqrL/esDmR72tVIRp+XJo4KHrgfQFsQRqUkqhKT9jmehPK2SsrMaNcHr
ekjmTTKTUte5Te7yydSwSBBGRjVaLbOIz4dfd0sRLKYj86o7yDfmGoRNf5NMPtFvMFc7wA/TMEUM
g5VfovXlvuP4f0z8A1qH9JdSm4uMQ69j9Xns3gcmEzvCC5AZ2dNYXbMyM8iORIqdgCAhLuzFmXsH
fAtfsiNl7q2RdQ8d3iJ4Vb1FbpjrL8jQ71+g5sZM6f6HkL9v5YuJ+34/KIJDfWdSbvKVod7l6qOZ
24RHbFC9kyQkyim5tBkb+hvYe76Ish7rOt3VuQqRmEpsk3KXh9UYEC0JKZF/0JTKearnPZwtZxEY
APsCknlmgq2uNLMZ75x7S0vcqSD3JvIi42W7UytUO8Hk5VKtXMVwLvBcjrtH0tHRZSSp57T9fvmP
PcNCRlA9NQV5w/syOP9ca31YmFUffAwbe/FtvqcgBNyqkHOM/QdE7fhfF83s0UJhgXW5fM8XUtJV
QT3w4K8axFuSnX+qi8m4gu+D68XHu5IKR7vWNtLoa+k5xb+eFKxfau459clsKhx2w5S+4FGAENpL
7+U2FsvUR2z3pZDjlcZpfwhkHI+fxUXyPS096iMoWPkifKSC5+1gifTcTX2LFw8GsH8UeNn80N9d
RrrUXaz8tnYu79AWzwAEvOudX3EmEsFM5Wdy+2K9lPNJATsYBPXC0+uvh1oD45UqdH7wWXEpmE44
oI5+fHkvDdYzFJje2dPFWRjj5uUUNLbxpm8ddVGSC4LUEGPjdEwUav18TKrC0uMQzNXBvc/BQTSw
si+v8+ij7UghUFBEig45tJXWV75GPNojzxN+ADleYpIp4ngWxDc82k0I05nbvUgdi3pbft/OW+Qk
M2Ee2OBNmqq6moIatzHxfwEqhRiDEz5vTYw6xcKkNiRxR1YR+CxT1/fKRrAxHtGfWajLjVNtI/Y6
DvTgFrBmGxKt0yLDscshGMjQ2Btgq5opNvCy/bwXsHqKGyWskRX0s1wNGyMgn5aXQ3UlSvrne26R
EryxV8qLDeEsGCLuyUANBNsZQs7HAO7Hpq200jotEL3BbyBIZPIFMvxyX1lqKnTmJeZsJj699/Z/
PFyypsFg659TNjEb8bagBdxLRZkpeTlOocqUrMHuV9i+f88nqImuyHnRoRDGOHgfMRKqFvPeVGoO
Bdc7uj0MBb6usV6vxQuOnHqyQf+zzbJxZoqRl0hc1b6DrPz7xD5ZSxefteQBK7dxkRZb5l1lDr/g
L4Y4WlEU6JAtdkOUETN14T9VyQch/iL0QN8Dnrb+fAvgEzPz59mTNqt+Sa2cV5F6VQ684/l4AvwP
Lvrldzjuhku8XujMZXkDDKrWoE55+XZanLwEXmOf3mjn2E+2m2WdVlryKLbCjaiVvJkk6EW2VdDK
ojOR0wjLgg6o0e3aru6xbTTMr73s4S6Rdpbj2qYM6WxjRqDBMfS1o+lVOxAnwIKjQbzL+WxY2Rg+
a2Y1RpJznxNSx+pr8Rg6tnHiSfPzR+s/3K5NAvh5jhZL+pNF+74Ag7dpGl6R3aBlHz8SOB3Nmgsy
h8Bz2J68Vra4fQTMNpT8JB+xfwFVZlUl0wQODCxEWLTK+d8uci+3heBeFvmG5YGRjd1zUfvWzOUt
0gQQETOR8JiV9MRLEDTRtE8tKE5xvovaGP1sB5S71do0z1dTUkW7XdPkQY7E4OZZXon1wweRQeG4
PJmr0/rZJ4GpCQTJW8d5hMt21qNwmZMJOUL99h1W6+merKrkISPl9v8VSzeqHmX5wztubYjczsA9
7PNo6z8juui7yU+xv1yaXN+HCnInNwQZDB/tX5i3902WX4sBlRWYKPnf8OaPtp7nrr4FRuax/0zh
yztfyaV2BvwibawD45T/a991rhTJdJcYKIuHCaJrFpJWJV+7nQ9JsodrIIw9IuTowJLr6n1AIcK+
8jAp/vtLNsXuShlYOM3mtDoqDlf+6GHEtl6dbPHKlYFJQQ5lbXL7ZN3AqTM3Eft38fPlBWPkZTkT
5Q2+zeTbw/d6BCJLelg6waEQhRIlSwnWfLJtGGUfS7EJ9gSAGv5Z8BeA7JqLZqiyKyv0MkIRTnyN
IfhZWJuqqQ6xeZvd2Hf/rrvverxjzhmyJgbT1vUOYcc3bwZyhLhDLPSwLjVe8IQChyMC8N4EfRu1
+emOC3Wj/q6/0K/E4XfvptFW2HmooSyQRLjkyaf52jIMThS+SdsHjRQ1QA9FYP/xh9+tnT+opI/6
9QmWFOC/fyyGWPydKev/FCM3ify3dH6QA3Q2bh2ts8sA2ShI/Y0tgoIpFpYS0kUQ5BwFBVgAw/ic
g+rhvpZmfgFAYoMu/ovVrvdziQ8QkKe05foXohv65KBVmJTCk6itQrxlE02R4cjTb/sZ2LkAqinw
F7GPF3pOPCdF7GIAyhrS1zE6Gishxt5s4BtpTxGMiLbdoe/Q1ujy8iFMFPWUcXMWHrS9azbOfRTq
74BPiCRpnr35/JwH+pPcbR2u9Vd45SCWclLw+P7CpHXBiCEbgJ/5e2OjMaqflmf7/ZKJacZmjsMQ
0m0Z8NBZhVOg0gaT8tvlhxOXerQ1XrCkEHY57dGe/YjvFjVqYK09BceHO5mW+ADgTqxQlupyxPDe
udRwbI29+7ivfx/UpeQ9cuiGIhz5KOlMttIhIk2OFn2pHv4u7q7jqdHj3xa44Ykp4/yIcS2ExKJW
XvOI02YT6CkIhjxgc+LmgJtdxFPEUcW3DqANod/vRlpDJV5p5QA47Ho9Tz3e3UPZS7wgoOvYY0VY
rrAuSMzGwpb4P99kO4+WdY6G55J6Ihna/TirFgXfv0dV/1WAi6hax8/w1Sn85F9A15f5vLqnKoWm
eZX3hSR5JCp0zOK522qqHMqdKIfKC9ecdn/S8e0E4VziuwZzgO1fCs6hZGPvklW2w7exxMur5172
n19oHixHKtM+VO9/J0K1tD+Qxw5bwQSsbvybUViVCk8keT+lCbNcv6WZ28kZV99SskNh9bgQo+az
4SpWEwRxMSWOYd+tSm0mFhfAZxKrcqdf/9ot04v7WXfYhvDCXI8eALutSWjdsujFlqdOxXTVaeBA
lV1eq1t7DQRjJvgSd2UJSFXo8q0VQpbLOshwH/e5I2icY1GRK1zFNlqG0mNbFLNOdZ42ZhcvXqxd
32aeEjIL/OZaoBtpE94nQcrtbbInoCFdnxweNKOOL/YGSUUXVdxq/aH2/DkoLl2ojB2Jothh+NIt
jGVt3YhB3le7z+o0d7GX5xcZATL88S947rIXhCKDIXhLGOJ86SYdpsJznlKC6DibKJ0Gv7UI8Hm/
3tANP/nVRw71kiJ/E/772DE/9DGVLfQ3MwfhUPCmME632W0m4REFaIMXf+u7xNUCj+njFWFpdiK+
yv9uN2ChXaNjac8v5So7dT7UyjMBEfv0ss9mAKHzy6U+uJ6UH7ovRwO5eZL17a7tXZWPAfvPrBVZ
GWulkywnTMuMc2sP8zQuCWapqxYom8vdJihPNFLHFDCxpowfZaGMDNZ37TjKPG310xVnDwiqsrvW
HuQE96SFIvcOTsUR/slW70Q6mneRJT6QfV1/4cpFRFEJSOur9bKXsml5PF18BSj1SR64cdnv/dO8
awYlc8ADH+Mx8eqpiYiLl3q1zc+37LOsmKLOA4dkFzWpbwCmGMjn+INhRB/Mm5kMmk1bSYCHp19F
ZXti4bhYvWw+Dr2kK9t7k4w0okvIW7x/A6pylYmpNu0xMtFcaGS161qE8qc5qaKXjg/yT1NsKBGu
Oq9zSWkM9k8GVFP02KtBbAaLTNd2v8o32Tvg/HJ4VwEnlgcJmEmvZQGqSKfBzA2bN1PqYDhWEuoH
2hGMW9JDYHQPiklBcKmVbxBSWJS+vVXjyd29jY2YnY8443bWzM6t3dUYV43eeU5VPTTCSyJPb022
SVbHHT9ynYJP3hDXxxexIQUbdKhcilcHHzN6IcIimINcut0hmkeIKgsX9EytwklKhQjkmufD2e/x
67wtdgs3GG16ZJL8OE/gU0ykCkiVLAjvD6vbsLFjKJJzE5vvNqlz3sswPgGV4XmLy2jOiITf7JoT
6tuTmuaesYNn/yt4HnK4g+GRzryIP+UnkU+oXMn9Km8zzjF95pCgM1yAn8xwBap13mEyUXqjAYbI
1VO5JPUd0igKV8cLGc76eJseat18RLU6jRblP/NtZLjgTqV1Gywn/qM5hYDVCysm0fYtLJUFsEk6
I/9Z+JP3LSUBVckNGIDJWDcnzeq6I29ZzMiPj+DEn9FGeoxedhD1CWpK079ulDRfjKUpBNBCCKM3
r2TD7OLOxXoIpPyLC+KsQimRYOO8+MjQJ87qvkD0SdM/d5+usRAGNuV5FQmxXceagGGR+LutL5U9
Dtp95oLUPtDTSSgF3LNNFtFI2p8tz8EJzzF/Iu57reKrvuZuE08hXBbLhq5DEo2uKEXHBAMePFgV
Vsww1F7Cg7h6R/08BYZ7hPaStiyt2wzxfqvNv/qrYHW0H2avk1SWoRo1dR2Vdmp+frkFwToeQRwH
4gesTDqhMP6cfylD4bw7DgUgRDDBBgtSP2TRmXVC7zvcJ62vDVSIxrbaYERP7Tg6dLsYvP3bGjtm
CscwbeGv57CIkEUaucEwpJA8qs2XaD0ADuUoFO7Ok9HGUTyfEFkxrbkmWnDjpGXRn8qQhc4gbIM0
pCnTJUaQ6XYDCGq/KgYxJTUJe1hwc6HZ9P/Ye8R35Idp1vJ0HF9gJxost+E+ryrIDjnzxx40S5pB
gCm7412W5+BqOdHkdgdWqmvXmYeESxoINTHa7DP7kxoKz/qlqPeuiQa2nkARj8jDiWPeUezSwnrK
gHXMN/Ne4AHKZtBT+Vm+/yRXg+j00p7q/dfHovvWSKDHBNjX0J6EL7x4gj4ge/Bk0TufaYMunsHV
yvGgJ0BxRk7vY0lC0tKuyXOnSeKbol3Adx35xKeSp+3VqHe0rBpJYkuLRKoP613ORhIbSdoLgLwO
64EvIaUSCOtO9XKinrRxdtQ4EvWq1IsutaYOzvEIdTG9DVwW09lU+o2lXUhhPJhrAP0JV8gT2SsZ
R0kJ+dgyoWXmSuHAHBxnf0tryysn4ViXBEMtF/DyvSKyxloOs5MUaiw7eQ673bOjbxAYlfqeiJai
2gtkJKM/C57toZeVmVjZK9SUYNaFnbFixw2sQCuEH3kbjrPhBr5fJVqdITBJMQFAw/ubpJOz4KTZ
LtX4m5VVmh/k3zsoFVvWfHIGId5jM0LzdNpmsKJlSw0I6th3bseGvXIyH5PevDeKO96x9WzYWTRu
B4NkcMA+jKXHeIxmNn/jpcjC3AHC7q8zvhr0dNaRe+EUCQYn2clUUQ+BMce2xBz5nCGC89aDEEIo
ahkyd3NIt8aPF03FyS8UxojrxB9+gLcplZSig8aoQWvkKDbBQ5irDifmcTAdhSK2aZx/QlqJcu0F
YcjAuQuJEL87gWNdBAMCA1Z1xJTe3kKsuymo7hhjennPf4MRLbgC2f4sVhFfmFU8fDDdRVMCctKL
2Kqau2kLCC9B/WnVHMQliim4q3azxefNfyq9mCCYetarhZjfyOB3TLb0IPmtAGHeClzJdGs5MyR9
+cfvbGSrts8yHtzOM6tDwVAN9EeM9zrMXbs3ULOUazL0+SlGAm0PIr+1p2mHyfuoxYp7e9dqgD1A
5+EmukFW4YPq/97UrIbog27ppZ3TwucG1HXVX8jC9OKHMPeVNu67h3xBgkVy7QVPuyBq6ItRjJMD
dwPmIwT/DD7yvpS6hAZRWQeGGEfintTAWzhiKxHBwo0/dLm6165AHhdTAdbFfUgwXU39q++SNM+d
3ziYdfI2rzxUmsDgflKon7DybsfEfv6Mc7hZDGLCS5wOmARCFuHt0LlIDP2E9k0aKt7Ib6XMQ9AN
DyTEDBtwhUlZ5yGPWJnqNUw6iSlEFcmzan7SVCndMbYY+PRH6gTlNqHexlewu/WJZ90e4hZAb54A
uhFpmb0htRn1BQtMUpIhSjPC+OOExHJX4J+Tb5dqJUyKOuTA0x+EmrsQvK0uRTvXW8fY3rv92HbG
/O1x4uBeqWA4PxlYrSB3xoDV4w+OfVy1yXV7vNa//BYX00VQ+K9WOTkeS6+hROrX1SdcOIKgXrSD
z7OJzEkjLVrErXFq3P26x6POZBQODpq30HniUYidD/c73VC0Bjp4jpaBN2t/CsFgqJwfnKDDBZyI
HiikXL0M4tYpNwVR8L4au/+kasrEcl8bs0tVJ7kYN6QyPjkq+mRLD3K458o/y1uiT/cfrYAbHH+G
cZGnGxqmkRJ18e/BZ97ZGllnsZav0bFSeq03o4JMCQqQ2FNSN++n7UeZSHrJIgyaY30e1PC2Qjj/
2di2B2rmjAZFGrtlkYLdpLHkFhf776ENZa03iNGa6U/xPWVDrjvezvjs9aGr84Gm2dLxLD+F8ftP
ztZfz5WPt1+I5ms+RxnWdDQq10NoOA4wT2BW9QnMdjXk23gZp/CryrMl8fy+JwkposC3S4McbSB+
V5fXLFY62YwxeiNiioV8kigKYWwQYDtg+p8w4VFPnqtsXkFzWfs3sxNDxnqfuYNUGWvKxf4zuFyv
pkwEG1/nqSkdUFHm3Bi1oLUN4yUUZj74faTaI43HN1yuP+33FQ3dd7yMn+dNLtyhFp77htHfZ25W
l0ILcwLfwKwbOWMK61YtGrGDkZNGChWLNZJ2WZEBQm3FI68iMNoaTACl19ID1nLd+Zu4MI0Wvdtp
XHok3adVMmFOGLQbyQZXDQSpDHnqPvLFbKamKJLbVTnp35i1Hf2ZGr1zRAmfZ3reVtmrKQTkMYyG
8MliB56lzhbxekJMajK/TtPKoA/9ZGN8Pn+2Tb1VJWhz0YYOT76IDcANSziOnCOio+qaL4kpa7/g
1rgwyHQhvrj2rI+/HYD0LFSMMT9ZsIhSOpvjKkj/BbgyEI7R3hnejrs/TXTqrMUlk4KW9vBOiBWq
1TxIJyEDxMrigNwsq90bor/L0jLiiS3Y1kP+viSd22k8v9goUlCAwPCw9Rwpv3/ybEXkRFAfjrAj
iB6F+1Nq62AM/JZT+a87ojvmQfufBKwz3FMjbQe+654CqEx75wVZKFdjXxUoHjzYf9drUN9sTsDj
HVjWf72pxBt28ShBDSiDOGK7TTVMRvHXBvkzN5SIsHaJMFFkNqQl4mG4AifIVqCs9gYQM+2EvWdG
SoUslwnfPe/m/65QDFqZM50rafjL71z20ruSRNS64kZArwhng0mLKqUF3K8goW2H4oVKCX+ziGIO
m/PxNKx7sNxYyTJaQznrbj3Lh4g+NCh6+0LrZke7AYFDUbWwXDK8CteYVoX/dePZxj34aH2mbhMR
U6A14sljHUvA5GVfYNXH0jNDZnqXh2miXRcTXb5xJnhINS1xV5B9JaSkAgn4W2chT4LsvvB/3HOk
E6Fa32nO0AkviVfZxNHQnvv0VABo0XGFUmxopZiQVOBh+azaBryN4otrQ/kdPycI6QCBpJETGyDa
6MyEpe4cd73SVg2BjMK1VIWzij6n7D2X49lnMIrfMb9+KaSet/0pN9TUZqJBDsK4OpRUH57FynR8
nRIZPxyEIoOSgb/mJnSKvmCXrxINczjmiXM0kniXUwybVfdHax3EQjpokCSVEHXInf6qGC0pYjVL
K3o1AM7J8W1n5fPEpOCx20wbQO/l3FDz6PIXgVQU2fSywy6jcW6VP3D7wwHGmhqNTY3pSImnNGRF
WHCeo/BSo3/u1VV4/czT68alTLysDfvItEsyYYN4iKHTSwzA/Q5zam+rFHTBJkFc2I8XVaNunSEr
M40IXb14Vbvs7xq4qwUpSBcHP3kIO6ZI1DyHnLsZMfP0gng4XfgQ6c+6K+hhpUvcA5Bl/zdhueZf
HeVeujwjdFvgzoJJkBTEuAbPkSUAixxHvxOIgf5Eh8123XWBmBu6vYTaw1L3H6dsDqyXixqsIwpL
ymU6CHhLxrYF3wwZzXEVgE/1wEQXkP2MyylOrfN4fZd2Dhc0tzKjCwxdugsW1W9DYVZNPoUuDb7I
UKcRgVQ0MNZEhsrVPLGTUywTHO0ezsSyXWrN/+DvDjcbqZanzzyznnTypCuHhy9JiDvi1zOwW++L
QkZEObGNXEZ8tQZA9CuZOq4l4RP2ykpJNfiWaZv02zqUss9Lm3b663tD3534r3s63i7tKGxedaEF
TKmCi16V9MEQqfLDnqT558euwwWnYf6hG37g/E5fUB8nRGSlTfZZmgbf5j9aeKrZQIqBnbW2eRen
hxax3ehXtuKEmtR5xqbClAvg8xW9Q+2x38KHFBb0m+ZTlSU0fgYQ0GClKXQQS3dwuK8zWpIQexcy
Un6ulNtuCn7K4z4I47Vbwd2TkbJHC4qo3dzyymxHjydJink1olfSN3Mu0VrdgLlONE0Q+e+A+E+J
khir/T/y43/vlYCLgq8R/vbeSRf9UoCxzcifhhdCo9rej5EU9DznPpmwnj1tuHGXqlVPgeiEgLrJ
gLglY/Sx7LeSrrwoN+NICqZlyTd51HdOo3jWVQe/cN/iV7k4f5eoguMgF0F9euOMzAwRSmjq+s4l
tc9q4c9LXJxREyhrMkwVQjAdr1n/sRThBfwcXgREf/pt5Q8G7+MX6nzG3jkChtl4YdEzZTXX5WDR
OFt5ZuyzeZvAvyyV+qNrVU5nP3zYTxToXXNmZcY+R+qiCYjp64KJwwH6nQd2fmCXeqEWcx683Gzk
fzG6iXjItmUuYJyAFg+QmiYuX1opaYwUGek32kaeHitlnvIs7YgX240iWrrm11xjBKOpq4ErXUDs
mXOsJva+T7np15SH7LJ5zKeb+BDiA1FoalgLif/9/MBj+pTpjFugAiAV3u0jlwKncdRvybkkRMAf
1H/rgiVyOj6V3xPHPmI96lSp4/l7vp0Oq0t2GUHPUTdbUNMHqee5clGen2KelpLm0DB2bv1BZSH3
lNHvWKtyQkChWounmhIJsMTbqAiZHJKAkaQbylBP9/M8tylF1D+mlzlK7dmQ5XdNxOxUJx643RN4
N6DtdSZChGP5D4n5YbOOI3bXL/xpL4Lxms3lk1oYCE1UTmkC9vN7tQNaJ0O9cfAlAp4RepW4uAHG
Vk+UPAWQss+joeymuZVgEJBZg4auBcP+j8GtFeXluwT0l3LL25i8bpuyY6+YdF/+MEOcpNWCNa+Y
O+B1qp7bVBKFV22YkaWwy+sTRijE/mskpcmRLsf/tvkr76zh/SiaoWg14Sghglh9emuZfMY4aND3
yS5Z4RQxZ2Hx0fd75791XuuSsYygHmg1CjwmfkCT6Y5jpB+WgR0QOYKgFcxDGrA6zI/DiM/M7KDG
/rrYNq3+0fUEe3nDIbAQr4yf6E4MFdWFu9ec9fLf5t4XgJ9NFVlEp4ORNKbHDMkShn8L4UTNwn6P
5RLeRi4RpG3zj3b1ncno14nqvQxiyxKpP7FOPF3KfNQgvbwkcScK310hO46pN2+MWT20JIZy6woG
ivyX2YA31wL3tGl4lErxdAZ/NAay6McNyAkvtvQ5dLUr3HSalTjVYU4vsZt4AyboOP6Tu9pipMzK
Ry2ZOaKg/HMKvZexI7kEFJBVdmWR4SYi06e2KaExTOaqP2PQer9CQdUAph6ipdEV7it3orpWwjvM
zmJAbfqO7xjShVyii49/5yFRjfCXHynPA5SFjZ5rKnhSk9d2PrIl6jCAwa/zZV+bI1rJubVdnAdC
UfEOeLULoWb4kvVfR1Dl/oGt/lfFsF8//oSdhK2BWK0SrcyQBw9ZJAdAWvQiM1PMr/mtBcNFuqI4
roWpE80qNqBd+nJgvOlVsKJ1T8XLPMm7tsLHw270xnJ4VJzL+VuOreCqSSgl7mTQ10suQUJSOIqr
ToaasexUYtbul6HSF4ckkZo30XVG3sWBDS2RrGsFWkVPF4ec53q5+FNja8BSgZCGnnV3u8jS9kEO
oy2ryvI2ACTeMhC/nOjcozgtqJn8cR8zE94ZlUHvw2v9KlA57ZGBmyRhwJgPWwsqiU7PgmZEOh52
wkz7AEVfMadin4sj/aDW+rX/EMK18ZPUZY7HfjnKwdWd7uFLmpfgbjxb748676gF9aY5StNsSEeG
jtcyIexFGFF3CjGtJfkwjgi8gachkfnx2qtM06RnDMaAwMJS2IRdBp9YREJRBXVezXfX0w+tHYeT
PlIkjhZFg+Qr2xZ1+8MOT2QeRVNZqjDBSiP8nW91qBywatupsvroFfQ5De0vFYAqBsav8GfnCKHT
OqbxaaYTOGd0a3nrGZkbs2URbvHqm3ru15LzJ1XJ8j0nHyXW7KNGPcEBjOhCZ5jFv7ZW5Tji//90
YrbcKbjCdlw3m5BupgARS6MCsLs2ik0X7n8FtlEofS3OEpXW2IgSpmzDFs79tp2+XdJly9OaaRfC
wWvKe5DGDUR2XWMVFNFvFBQJwzc283rmwA8aWMYn0yQnNfJr57pcULocIy396A78EIHBsadLEAzS
GUfauUNd/ZS2eb0hGDTJ/E15Z7mKv6gBwihM2IL5CQORB+/rVsdGxnSIMnBfiolEL9wxeNwbUz2/
3wQvkMleYsy3FJTuK8NLcImXeux6rTk2nh5mcDqhPApXf2QkQcW9lz1RvEf/WJV9a/v/KKvWeSoQ
147EqPLizs7zOlQ3jO/VT+bgEBg/Gf8lUqZn6E/vJjuD/Bc8BPMpbb53g8ZKekwuzmo/NAamc6Zu
YoN86BtY6DLIWgWRLlBznFX9ITsHFTnjLmTwfg3XeA302ZxIRvgSGKd1XUM6Q29RUGqCn7V/wbAJ
3R6QbTYznnjZ2WYyR77ghKvhvie8DNeKyvXkgc/9bJ5Hi7QdLKQdC5oEFlg60Ezza/0dBNRjF24S
W5B7hhPOoCIlwLYbNTaR3Ps1yzTsyK5IVG8ysnmciEJRKuhGw0RRI4fxBZdEM01FsCscu8XkfBCU
eXoZDICTMp5GezPqONwo/auv5jkrJZ2TzEjm2eiMyQHBQczseYy/HIJYPsoA2SiJ4rafy4xNhkLi
r06MkSinqlvCxhnVjYVnxzpc159jCLNTVAc23uKUpL4vlnEjC4ACQCj/nJyRSvLR0TO/CpI2+tvL
nnIqwued/Do4DQsdaE3QZDVwaZC6afc+QWZMdU0ZfxbamH8NDhG5Cy0zbkkzyZYNlfcMpMQoDqxK
JMkgTvagWc3FgicLRSExviZ8XTvWKWCKy0vxaJ9RjMzO03uy3igZ9j63e02LnYN2Lco9yKQpfvh3
0gv6U0m2NGnFVeXuQQ2PTNyOsAQvu7xnAdppD4lwmkNV40QlH8FkqggjmVcZL5zVm8EMRqwZydY3
f4QGAkvwfd6DC+8wEewmRd2YRwtOM9s/DvjeeH1un9lNWM9wtyylYtVylT7/SISke554MoHpqh2Z
Uz3ORfg/QKmwUAgXtWgEHpM3a2imDI1jRDDQYKYTqr+QM4tZ4iKbaSAvdeaIfFJB+3z/63LLakIn
JeycBf/XMTPtYWCOOa9OxwijJl4xe9Qxj0AaSRlqDdxsL2eugR0zLnOvJujtOd/acu88NbrBZedV
lNfQtXD8hgZK6GxteVGMkLziAUmwaoVUpUYExOU/8CPvJgmI4HIp6CE6zS5PWLM7U8MtX+UIsrSS
0evmaE6iDMJ64yx1h5IaRiix+wx0T3CbpTYNLS3NIsLzCdZZP/EKUcaB+JcwpA8GTjVqT6rk0saL
gv2aZbM0sXCPCRZxuaAAOfpiBifiTYn5GAGJfyQ3Gu/79e4mtLZGkxx61VhdS4YYy5laDvENY4BV
rfmTygZh+uEQEEQmIzerHuVpUQKdymxb152hJe9bHjxByQWmEYmVcCZWGEUNxi7hPI8fgn++uXje
vZvOkfNVaVGqx33Yg7LWjKDcBKKf7/RBsKRWr4Zl/WFnvUahqwI7ucYlqJ7PDDNOVB9pzj6O7Sct
sz9QXgsNXI1e4cdbY2nRhgzT8VuHbWnZWvx9F61qwRddNbQOLmDUcbRm23fSypzzt4phhOQ8QDy1
6/mAQVD1gCiPk+8vUH073Oa5zkRpxcJcIlJ/7WNfC6I4TSJwg6z3OG3CvbZQhcdenN8UhtO0JFN1
vQdEKBnM2WppQwNwcTQzmFrH7CpfQi6eqLb+80XBeJhA6yatzSZzXe0HRdjXLsbQNTPO6A6UXDkv
uSNNEgV1Oc22Hghy1JKwv9zRxUR/BvLVYqeGH7F5TVJpRW4n8CfEy2hkCJ/92aJ2yxxMoj76hNbE
uG3ktYQ9YTHOyfFbBftcSX5vf5e6W4JQHvNwQbjowu/H1qONj57bu3t5BagRcENvAwBCi1lOtWM/
1dXJb4Z7p7iVu8FRIcC495F2NsWQEU8fRJGEdY0cc+ktIGrokBXGgrEKf0g/xWz2KVap8fhXyKVo
Gu2iCiPA5b5GtB7u5m6chhpCMeNJDNGx3rCN4bGbnlAQZp0RIOqhtLhU/zapACQt2HHPmumws7M7
X+92j7Y5BxGkeIN+tEvAjK84j3D89q+726h3jFKP0c+wQ1CDd0YHK2eYlOtQRlnTzM6elBbxiN3b
QfAs9AFPJiPtepoR30g2bK5PpB7+XX7H7s2bHEXivA7SUDzw/62qpBUTsgGcCeVdOx5yzdP+c+Dq
P2YcHPWjiIlN3HtUzUZvg8BY3aZBxkkrYFmCpELXSyPYR9xl3TgEzdzainaGKXfD6fS4rgtNQsLs
fwHujuClflXdXW0MN+W3rH7iOB5GiZ5lbqegeG7T5QyihVBTnq4tfWe0mQfIyebpatzgBlFeNYGo
eR2jY8G6NsUXn4E19N2flqw/bzguL4oFz+pSq70InYX1bnvc/KXNSiBzPxdAbn0FIzGa9cpuB7dN
/Zdauaux2YJu9p1jZ19ZbTq/kkedxAYaRZPUz4bFWXTUOpYpJgC6HGqhZ3WjOBrwllTx+nFAA2rC
pYVL2e+kf8XM6zTqushvDwTMlqn48vw3gS6ba2ctuR/DR6pjQX7Zlo4i8c+KKYROdsMzuBo+eSWr
088KT0z/MkdE1Zq0HubOcedUvcNLsAkO4AudZ51b+h/uD29M2zItIelsGSUxgfF0I6bCRX/Pb9Th
6Dt6wVJZTgaJBDWMTMCWT9bNzxy8YR+lhtkULArQfmpL/SFi5Owmem71LDqphsnNIaXpu9dsSbsf
0FTyvpPEOannlB8ydGL0jTsMNhf4u7ge1RFfIGCvfEj+apxd/u1bk3h8C1l6pCoOJsoi+PgbEZ7y
c6Zus+InEDCClwiFVpyLxVXF6YGXs8KM8qdSXTTdAMg10RkfBekYELxkC+vGejpGEVIHWLKNz0ny
vMCKVUcYFFKJyaQaJEaxhaLNs2W5LjgzOL9fxMilWM2PBR5vsgTugJHETPeRGmUPXgsMG2xIf5N1
9D/QgFu3Pv+/eHGDkhDOTBzI/su7jo6wUI+3VEAIGdxSANQhIGna4m14rll4VFI5i6ks5S68GtY5
ttMIhXG7AeJELK3ejAkJm5rQxGQCX+cnm1kQrSW5KKkDTo3ZuL600iwrFl9WA62g8e1sm5Z6YLqO
jeUrgyDOghDru21fOZ62kDJEPpIXZDmnYRSENuo3PPJutrP3+QP/G+6rEn7Lzqh2IDS8li5AzNwY
7+EIX1Hs9arlDEoYTd5aua5WYaytwPxsNGMH/CCzxPAAz85kHcztiRp2C7Zw1QPG/F+equP49Zmo
PAe0eko6stDq9RvkszqIbueCWumvVB0QSdwzikeplnjklQ89SdcPXrrlz+0Lso8mKgkuRRU/u/MD
OjZ6mCJKdGRbw1eUUGj9rDowi8qolQ92S9Ri7cWEKPBQtWttcLdk2Ke297FSUSrSAdZIW/TUZrsb
Ta3LG6iLiObizV3FptS/R0/aPASNRwbqk1zwHtYL3Zu7/szoVeA2VNxDEMyDIk+6h1XRDjHFioYN
quWiqq88OFcYTTw7NPDz6Ktmwq/B5aUF6WSO4iJUFWAlE/It2d8E8IptT51B7ORks7xuWONyMMzB
0+RJf/TAMV2R+vLf6hw+Ax5t9iuyZQaHoTMwrSAhlCfAURDscybFGq20ZyV4WybzWwW21cuhZ/az
SaQh75nPtkpn9Ty3NZffQEi9VAYUmGNQiAhJitUMakNVn4NGLAP6CnMFLWeyVGifMw4ITG6ZLSEA
OKhWd7fzp5OlrliWWi2FG1fXyo1OA4/XFhzFRhxYZWBdAkHbZPKAM3vJS6KB5PnJ1MyMZ41/JLOH
sV/UWMmHcXKzbG/xV0KK6IfbPiW9wTT04s86xCg1LuOPhDFlrBwyoNS2GK05cXQEP5uCQ9pGfsh1
50A7dnLD6mJFyb7hz3UppIMYsqCmgY78RkVhDEpIj5YP7WelREmW1uLKzmKQVLLFcOAIZyfbz7ct
mWcsTfSlmWtiC0owvsqPkfb99kxDE07SHBIrBiwhhg8SosXaXKM4vN/S1re5SN+iIsfIic64Z0qf
iOBMx7/AKLenXJ8FEZA3lSYO+K2M+vX2pI0UrvNusgYCc90e+XZHJsTpWw80HYA+tI+SOEfFQspw
KH56eHTykhUjyjY3C55vbtLVe5n2ekcneh6wK4LvuoagR452E3RTYOGA5lRk4NxkOaVC5oqHOBUM
8SMWx8ulhQIy5xPyTMNtmoGeiGqjfR60rAC4ei3QswfoE7ZD1tSyCr4zE3mqXrVkL4axy+V717a1
cTX7s5IpdFxpdeLUbykgNbtniDATae1Kt4QHMlOJbv/VeZ2LGZ7sZSudeQLig+lMhUzf9FNCCIc8
pwLnfAOnho+47cCh1YKW0I+ALo1Rym39ctKDE0zmeQuEkjTMB7QOLQCc2IZOd2wWSv1w7wmIWEQv
8ZnwcFwpgHp9PwXwYxq9gW/0JOD/b74SwUOrIRedGP1LqEmNAsdTYUSueD7x/uE0Nyos+1jmsbLB
L7nwYUjuo9BMM5/N8IRH7oRR0jye6DciEf7BvGWPI4QS8iRfVz1/hLA7MqaRj6UNMFB+ylIZT5Oc
QzVLbVXkONTWA/QmDVgSJzjLnMpC1Y0aY7Y/bTHKrDnIU6W4SmstdBFBqrF8hrTj3GGKMI33ErsQ
U4wkdxwq03oz5Pmtj2JT3fRWBaAjsDRJFPcJNPYE5g8/SIZL5BT4x0O92Dmfa9zmHfYL5JbMC3YD
V5UEWjvCpyLcr5ypOfKLsH40Ppab3xAafsTIs7iJiHkcf8tsfl1413ciVzkjctTMqJisMC+2j3G+
2YlA8l+Y2aM4VNbULDjnwfcmZfBtwY9ObuRCKlm0aoQyNx9ec8Ao27HIlFibQSlgpBzq/mg2hkzO
ISchi+s+HAYkwVR9VWhVTOdC4RgEc7LkUSns5sFwnhufjkuRKSQKSc7iLzKYaCDY2L2705PyrVHb
nBYwzsFMfn5JiouKqYtQmJqqHkCX5zsk7Q67AT9TzFkGhZe71sv3BOr8PIXZGevpXIALJOztlvNU
udZNvTgYb7izvr+875p3zRRCV87seByQz5rqikhOv2KR+Y08EGHulUBO17o8fbPkluUS9sBb6z6c
wx+m3AdVDMjy/ZYtI1uvqFjXPLoh3yW9JIr7yofoHF6KqHYoZfVNdrS9/1PEXGaD9QbLergY/r2v
1PNj9HSLVy0P84wxG2+/ayLpEnE+hL3v4xnAu7jAgTsJbzntMuq+vT9OCLvw/Uxxxc2c48iF3xAB
oUAlOcXrAEeBd3bRdFwci+9GCWKnYHZHeGu2mpBJZnC10kAIr7ixUef1L4cqdFcnvB8Fr9BY2FaA
sQGSNMrhA+ZhTKOyNnY8eNJSrhZ57cDtC11I8/Ltr/sgo9YpgU9S62LbAjrEvAMSXQX7cmRfA9nf
kd7kTn9rH8CwWgmY/HTX4J8CkqTfrl38ZdchMNAyPrp3OoZ0Cnu+Q4urbpj8zzPn56waPQ0YfGUn
w2QcQCYebCniTLkhZ1Cveu6n9rSsCI1SJUvWTMI7YeHLNmalWsy99VNZpDvPAcarxpYjRP+Csn3O
icI/C0JOz5sjvD72Oi6fey19obe/FSk1PnWn4HUnOcgrj2GGYzdLGK+n8nbDLN68X3Fy1qaeqjyP
KJeDQKNqztGU4LbFq2VL07ClOs/Ttpyep3eeilxnEl+4Yv8BAmRoQ14tBajCDAVPsQ/of/O59aLk
JbHf+Jtcw+rl/RErtSMDb+iBqflCzKi8KIx5s04gJX2cWxE446OZ3MhB2yUGjKZjtrMR9KUFUEIr
ER6VImtXznuT0r1JNhLlPmuPP4SJw7VkT8qZ8pYoMZ1fsX77xNPLMKG5RogCfW/QfcbyJdaK9j5k
z3gBQu7ciscysGhDAsMPOndopu7ZAGUcqNgX0fdk3LQlKD3OFx/89wjDNoxlsfInI8feoSzVgfWk
S0rE8NElToyH4fVyjrl0puB28N10ImjbWDjEct7MzYAaVbraSNKGpY72fpEboP/otaU1rPeI+EhB
KRPSnm+O8D661NafgCDREseo4avmbe3XOQHFZL6/jVidqNSra7hCSRWVoXs+Qs7vbwgR4nw3tpsm
BHQzf3IDfHi/guIWOYUhW8IJF8qVlIiK2wBEEEglhl9GD10V3rWXIc8sz0uzvQ4ULs9Q6n0Ridez
m6rzpoZNvsikgD28YAr5maFNiNqKUOXMmV9h6ETfW91azNXu+eZB5xA+rsOj4f1ZTDKUyrPgU0gv
PMdpEAwDihHWWNGyr9vyYTDsjawNRGSNo4UwJcWwDXy4/III6ABHQkq/zwb5kglthprBuBcE/373
pD+dxxQZkLvTDWAiQeGwzGLq69dG+yVgo8E8SWeh24TlNiZhZ9bV3UwUEIQVHgW/jZpduEJZKO7l
0T5QwY24MqXSDr0C+PqDJwzL/l5VswDwilXSESMBfcW8i+wrDOhRly7d7BRp2W59dd2qr3KyRrH+
3iiih2MP31t9jM5kj0CSXvhUknAIHi1Kf2xZbDOIzEYR5RCvpTqTXYJ1mmMvmJ4atbBRyUl8pkVg
We0U1KrdsW3V5tTEbwGMcOBGQ60jf+vxnKkTm1qLZo7lGlKEydEEAdszM73NVhk3As4LY+SeFcYc
MgL55gbI7X2GQsGLkK2ujZ1tn7AQLGXykX18SCWTTbT6u8XNOir/mBSivF2rng/oArrIZwqT0CKd
l827Mi5L0JOfxCht1alk1fi7Ee+tzeeudQoIcmwVKoOZRCdk7nE+GSmpTUzKH0HVUkrLXKO1qyli
pbL2KYs0JTfPI3eVpwCd8cHJMOQ9bQSOeZG1jkgd5w0/c9sNfrP3bwT/C9kB2bqKgn6xoiFn4KBB
mjnfS/oGQMSYr3PO4n+4/dW39pY1D+HZSqDhAUn7LJS1yudz6VFmIjvfGzBctCP6B7aaXzTH8jSc
opslUqhNObuf3smdPI6uyRcZ4xNlMFIGYYuolQJ9z0ch5guiIyKnLEGa0elXIAol76K5Rivi5ym/
evIwKyGpF+fEsysjWsF3Hy7zd6tQpKRzEcqCZ3XYD88HEJlHcdVZ3f47ZzgyHiOeO/39zoiaGMDk
VBEcaVjeN9OJBcQka++6LeIi1zZIxtmzDdK35FtU5rzHYv9EHzDPWtUOT5BLM2DZ+lfguPHQAxam
1AzZW8X0v0nMbylVFJNSxTZ0Z+/VDO/NbLvoYOqDfARitBLF9LTk8q3T3eeKmHg34Z7tdErg0G2H
tfyJtnKlzitYPlCFwpdEpmxeTkE2Pnqid2JwNGtL3SdbA9netnrjGnGL+VNGJKAFKtOruIg78rA9
CyMWF5COplKtUuJESrOQTiAD+ZMfydaNxdxWOS2mW5Nj/3H1ydSB4euQrYSJuWvKmCY2C+VBYOYj
5VzkGpJmmDcl9ZJkRT6qGZx+wyP/do/w5vYMsbQMTW1q7Q1vbA91lLMIUbC5wDT61zrk2WEIIAbs
NXDE3HCBuG9fSzRkqHuqz3Sg9riKw1Y9a0FrMaDz9d6kzZBA60MO7T7WqbaV4Tja9j2gWRZQw9AQ
jmOGggCGhAdf+WcQKY5o6U/9PRpHV3iVcfIgGlnqN9AoZ4zf1+PDeTW1093fP2G3hmuyB5wzpUne
5I/DTDavh+uqp/7GU1PizGqCzew7JMagMvSJyLibFPJoeDUu/K1AWSYF1Cu5ywZHoV3/JSewkQ2s
I6BVDHFqJ8R7G4zLvvnzaFe3pbkHVi5IIUIIcAXKnFJRwYKYXBswM0w16FgoMjSMiMfozqHVc2oY
5MaDZhFheHszkrSN5x+ve5WThK9OJjtD7wil/7rnF3VoWITdFVqdDjolZwp38bOcLjy7xaRN6IF1
3zw+Sfcg6tXzW0zkhZ8KrdeqZuQSpB4IZ8o0Zkpi9c5cEXDagDFEIvCJs8hlQYFxHZqZUi6GRssi
FrC9WfQcxq8udMERrQrIlLfbw/p7uvHv8A6G2dfneSChKSwlNaliSkZrckytnilbKp3evijW+3J0
ofp96LdblHS8KYj3X5bZTtah4yqWzFcxcF2SIk06+O1eP85g9WCaO7ErWxUuiR7/sIzNlidLa49d
3kOnfw+U6FtG4hK8d+u85Qv5YlhNzpf767Yp4xPBwTmy1tP/6SpwOKke0TIvgRc/a4J6EfYlQC4P
s90uRR1dcAk5ueec8HMf+lICGmW1cL0iQn0HoDTd7gTAcYpZu4+nu5R6VTM7ukaU53KIRtK7yaR9
LvDQT7pi66aKv10Vdn6P5EsWD7Apbgt1/xUz5vXqzvn+/g7rtubZ87JRWiObOGh4wIMsNQn/N2pw
tVIdrUGePLtmVFxN0KOToP+FOrVMSfdTiurXvsA1uPeI8AsovoV7bp+wjwgynBR7TFmDkL0OR4F9
aZPYGLxkWEcBDXT1J4l2kr96RRPb6ky/eo62XOtyR0J2n6Ro1iVZ0RS1423ZngggYHlBdSfqU6M3
RDSgleKEJmEY/IIn05QjVqC2HcEPXqajBOzP7FM60WRds3UlcrfsiH8gHCZqtus62VitCL48+k6+
/GGHzsc9MTmbDfWOgl5TBJS+VHPDPwZ8IMlcXgZJ5WWwqaauNnPxvI7F6QnR1BOTDid1AnV6WrF2
BBoaWhn5MoBV/B++HpL1/+G5J+x8KxQFIFmXj4uWaGex0c00kO8hvMMlPlUg9HofC/HjsX01I9+Y
Rkmly1jezUYaOvQYbKQJVMXJu6P1qpwJETYl/X9TgJ+wBNJTDUHbHevk/W5L6qU7N1LRNANtznnD
380n9dTYDS3EUFXI0TeH/Qv00Vu+f2KtQqVakBDADS4NOC/lS2+sh+Jp1bP0aVR/rLFdP1uL2hT9
eX20hTeTYARthBw1mTkKFZPg/HsDdh77rUbJ778iZXTXF8Nldx12U4PzbhxwLPCLoeGi6NqZjw2r
c2mmWFP/5Tz/QIRiucwbln8k3vwpt/3LzQFGH+lbziEUvi49GB5lRHe3gqMPc4nvnfcc/Fpew7U6
jUfkqzCRxfWv9WoO1Uy4NV46Qgim4r4F0jk+F49FhGsbc2Jlu8ZSBMaGfMZOwPWu8FFmBEyDkSJe
BtLqHEymVeTyhJWtbR9wlaVxpWLEodh1dfxfaIMEtpM8I4jMcP8pQdbivtpuwNSqHeqxjVh6kDge
QLydsfE3CxBfamn//LphmzfHdOAwqGgG77en96vevOcDylIz0iKbBcmWHX+o4pm1Edho9JxI72qy
nnr2esSLCQfgA6IE9DekI0J8RnE9I3aycyGMdv/ObqpDY9KXxaCb5XARZ1qAqMW3ovXEfdwC1mJ8
Gp8BFvT61z/mx8TWhVCyo+RK3qPw6nLdyJCF3/PyHSDv/6wce6JLJlbcztZFrPw5EV7lvybjMQly
1J0hsVAR3MaF2CgUxLxIpeh2orC3RlZjmc3XQLB/Q+zmEldm6YoMR+JoXhl69qeBKl7dXqUnsa1s
Me4uSdd7TRR5OHixH7o8J5RnmMwE4awVlJUFScbyHgrUEiL/e4Q6opryabgvLAJ8J5RREv3+Oopf
Tx883OgaBj30QFEIOAOPHOLaq1yj/ANbiYh2Csl2GbvrWbLsHHyimc07A9CmQ9BZ8jKv+5D24BQL
caCmIfjGVGC3xc6hcIQTcSu0dfy8uwSsocYvAxqk+kMOF4bRl32EHmdlSR1DiGG+DXPTM6s0OSmp
hq0g0VBbXH9Uy+cZhn7gAG5x6khSPpAihPdyaiqXlQztO1q3rHrL7brmn+t2MMpnKY5X3Op9fCiN
V64va8jWE0PFGEsGU4AJ8nLTT8ObYIvFRUVciTTHF80GipEjx/Wa9kva/jSB7+8zkfnp9CqjM9hq
Kc0P+vDOAmwHMjr5kfpMQLETzE+AGHsRoeT7/9UksPcumILkoI09O07oep7qZclfa6+RcKQ9CA+p
xrXeYsYxyy7T5+s832pvpVRXL6IJqAwsm8sm45WHoflrW1VkNx8w0sJJF2lVAQdqAtx7NA8HHLHu
do22daShInTCw1KzB+CwHt99chGRbWXYxPYE0lyj4IulNUZCwhI19ic55H1LfzdqfTbbdPWikHGb
9Gq/VgJh4HnmaHW4qnvR70wzlqFeW/JVpyVF/5kOInE7E7S914ApGIfStrvzkruCF613ly3Sn8z0
s4XlQqeUdN34Y/7eBPo0zrQpl5rTBEhwBakBLzUOn1kIs8wn0p+PwTelRL9PYW5EkqZup5HRZYHq
9Bt7B56RMqnOLUiysX0QnR8woAbyTN4kQwrs0JpnZ0AZ7fY/aNXcH/xp/YSL1WVprheYc6HbMuYl
CuiH2V48oQG0CmfHVMKFyS25lBp0SPqr6/U+yaCqFParBbDRZKKBLWxhHOnlwP8QdVscdi8VpJ1a
Wp28zwT1IGANnahd0cwzEYT/nwMy1hwtra76Nt2JJOGYCxKFyjyVVhiHjMVMh0OPaO65B3Qrajsg
2sGZJ12sZWPUpMbDJaLNL8sR4Q0Yo4lg5bpW8zvhUGGpCl4LGCOoGVefQppNdoQu/gqyuG05GDA4
5bnwHEdUM2eIVJvu/Fxe69TKJBn1Es8NS9NVCe8XqPh92g92D8CvZe/VILxG2uS50HncDwevUpuJ
ZXoGjxjieMZLSnpkgd1a+Kdjetmr6tffDXOt28cYbcJZrT2GTo5Qi6W1Ed2qhQOxroSRfpQOksXy
YJEzM7mq9FdVx7IuNY0OPbJp+X0WalvEoMDEC8DD7pReJogmlK2Df82xfxMnSyeaFBU+Wb0c9sok
sHCCk+D/BHTakPR0dJ8bAoSRN0ygaLcBZkHjnVpSa6sQaGBPK84FNEVzjCgOsv8NEq7k/fPJHpPd
vdjM1w9975D1rQa/RwaUi6WdFLdUPrRkz+lI0iZGRujq1E3cwu9syLBghNfDoF+pH0/J+diJb69/
VcbAMSYB7X/CiBFZtUyInDUYD9gk7cxnSXecRp6X9Zriv606gtUqLNtBWvmjhOJ+3CRUCuRuqhNk
z6ng4Ou7GLs/lipyePRrK+nuUhjvT1rVmN7UEz6N3lG86xA5OH5ew2boNn0ZtKHSayB9/gefvAJD
wNjSaLo0a8gjQ01Y9hNm6aCv70E+fgEf/5Ud7fgFvbV6twd0PgKw+UzndLJrapLLGXXFI5brVsW0
8mwnugKit7MJBaaOXmfquYjbRnqqSgm5+FtUb4a1LqXI111YAnmbyF0ND3XrZrp21EWYCHeqjQ+V
gco+RVn8GnVPYyyrAV2QPlerzgOWvfB5IDUbM8y2xsERoWawXhPbV7YNL/5orDHWSv5TVH6fr9w+
rk8C+Da3szIEJ+33h12UqmzkrHSDMC/Bjtzxvyn2d5xkosXs/pbJ1j9Emj3BPM7kfK1vsCTQ5fgL
H7xjwZTxtJwgpXjkREKg64Xi98fNUkUx6+q3i8siuXOyJ11Nj/P6b6prZpD3Co5wLLhLIz6XUNDx
Am7lOJiK06DZlx27AVC81uB9KWP08HUoihZ4xg6u/9d6xtMbF6xLIK6c0nBIYwu18Zmb1DmUfxPl
SCFGwBHADSRfb11hcpdoep4//P7lF+PiofjBErxwZzUYI9JJm0vjuqc/tTGFPGN40jRueUYpKSZb
IBbP1NGv2i3F/Y6KHVsgWE/bvTyNmq9fsxIN5NSy8Jes4zkXtjAe3qmZP19rHln0qkM5zFKPoSXG
MdgVMGUM7gjFsmdYwoNmGDyv+Dm+XDpv2UxIG6gqZ5CFr1/FuSIOdSB4zU9/sl9UG3rONzNbZuvH
4vaVN8WITMYtRY1sjp+Ox/bMXPOPIc6HSUs4bp95/Me/0nmDe4WWvVLRFS77/xqpI6LWWjRNdDOx
NTA1c5JZMGb5m+Atk8XEMimUB+0dQz8wzNlqkNi/XaKgWBNJtjO4VAbyzBhKxpsp6XRLY6p/ZPV0
O7Lu/n5Y4b0ffODdodYt1Y7I20SbY2uTt29TcIuJhIhf02bxBg8Yg6gGPvUdzXJ/CrxPx6Wb+4vF
RrPzvR7wT5V0mn9q6PJdLhCM1BaO/cy/rvEDUC90AoMQsDxZQZ9v4Jy4iBTbHDaeHe0IPBXWPr7e
xS8k8sbD0YXus5O15nHyvmiFVFjsXVvp8O3MJponsC8X9icLNZHi+rSql5o4GQ8rJEuoMxF3nRRb
GXYhYyaFS3rfS0pJqBRdcGXf9NgpmSfCDryfQ7jLAxue+7zCrf4L5KfkM5e2Gvr0lVqQ8dOw9imM
n1CtP3PH8I5d4MgB1L1kXuPIBfGb/1wlpD0SZLUq+zSseraqvjQ0SqZNa7b5O5nREL7RDAH40J9c
JcgdeyfKhAlX9hC3lVgG2lPTd5s+RkQNZcMwYtWAniA45JFhbGnPs7d64qcLZQbHc+YkdGUlFViN
d8JTBcnJabQNyTfKX1KWRpeLJJWKP+S/3PRYff2jgDzt/uYWg05HmeUAxZTjJa93YyeiIWM6e+9k
Qxv3KM3V0Za00tAdARxvFc7EbnQiYIzrS20FmeXxenIkzJ94YgYWVSazjK3J9vyeyFl4PbSNNGQi
qpD2CGPs67HZNfoZ/J0L37TU3SlKdC7zpPYnlSAWCtsPCFUuU/9UnO9vJJ0UiXAfMV9N0AwlmS5z
aVajMTstvzXsECCMAVrXoFAgWD7yuFkjFmemqlsy90aTENkffuOmtRruD4opZJyPlkuK8TPHBBC6
xKy0V8Nfg3xwkBLkQJI1nMF1Jxz6zb74xdNJNlRWyWBUTtcULL6wtKvIG1Jb7hrydBe9+4ej7WT4
kl1gKi207dIACnrPwaMt7npnTVQGg4234mJ2kV/sGfkVpppqqq011HCUKtno0skmd7vAQWKCC9g8
pOkTfEyFTebLDl8j58ZxV3yIPHeSPHN0gty/JH+pm7mtbz6qBe2eImVusk4EicY7v+S4O1heBU8o
dif2JjbJ8uM+waD4zrw7hFfm+EYozeyq52ZX2EBrfcECfErdkDaeTN9gzPRqxCkmLG+nqxWuiNPF
IDhB83EOaipEINTv99sJpwIwWuqHQOVMM7imCwd0cOJjbOTnI/sJZ95zfXGzGEQZx6A7YHHvocI5
ZpoxXOf2CqVuBJxi2BiOeSvbei9SS8E/WN3UpBEszv1/XH8Zr0JxgdprsnYc94rPpPtDzzAZKnrN
e3BFq6RpwRidJx6aPo7rofpoRa8xe6hkKaa1gjRe3fNhu0/pRwX+yL0vdSw3CZfK2sfpgfUsybBW
8iFosmRgzr5QH8A0vhqGgK3av+kMvg/crvbrsrnuq+/KbmqY99AZauPm0fl45vKAVZ8A/j8fePfv
9tl1vt+YfA7OzeLchqKeJMyv1zUWvmssRwGB7UH+Elc5mL/pvNxo6zmJO4jfGarXilVz82SQUdww
MSvqCVba1XirsFu/oGhc0d6ajpy441xpB4EwOOX4L7vTmWquyyGepQ1TB28rD6+M2RnlkG9Ug3tv
cNEkglNoQEd1S2DlmEg74zbAX8qs93DP3aq4GNJmI4GSB0QJfgg/2mo+YOfv0tmNcNjkIaPpLppv
mLYx4eiVBlksDTgDb1sS/piU4HA3ADWYSEValf5Q295PfKVugCXQTZ46taBfaWZI0PMXod+PZYpm
WBlZ/yzmaP4s+03hXcqAgK4G8ZLIKTB93OxMlCMHPE4emxhbbMIrNURlUnw+v8qJgFbf0ggXK2Bk
zxMZQZ0u0LjgQ8KduW0HeqJR7WvQDvAxX0YZl6AsaiXEcBtwtu3GH7uO4fxiKUev6+vsHR7E0E66
vWnCCBkrzJ+TTiw/tiJvkA9WCpEpNqkLgKIeWviF0n5G+ZwuiPG0b2m0EqHuxBTQwtunkSOrAuLb
f+A/qtgzqmgFhCetYC2uVWRXMGhEkOSL/jZOfF85qy/cnjO7UB8T/O4C6KQpxaf7ccfL5npc7aJS
O6f1X3Wg6LeBSp/e3ksSRTchDe90HiFb7GgOkoG5P4o6jSXnjBqoJ896yskOV3gAGPUVyaOqpqmH
eZ3rEjATZshUEMg0E3ZK4hshsT/fAGO+jx8xvR3Rbgm/v90hkoq6Hg/qA532r9pdWF6hEi/G9Rs1
my6cxepLj/7TCoTlk4D85gossAENkf5Q+vrpvUGin0LS0opxA4PvQbjYqzJTnumo0/4rlaj8j0hS
1tsOIxNfn6PB4/PSafqYCMFphL0XqXLQhbIwFF1Kzerqper/VCBNBphjdL/EeUoxVVaY5AaZp++a
oO8YE7PfLHRlaQ5Kl3MYEWO9rZ7goA0s2DxjD7jMX+pMuCLXQwFz4TJfkDf3n5MXLIRKuT7kpvvh
S7hzjGhu6hN4bEaLFK1FIeLVZcXCujNZCV1QSKNXuWVXR9Gkv+9LGfywEG8iLP/K+JEOrMdVf0UD
xCw+9J+EHj21LOSC6PIGK91nFTfkSFfvBXRc2jN/VK8Kzn8rf7/f/JV57+x3paVg0UMPmE7Q8c05
99dbOIDPgv4lVP1WxgHf3NMImY4PDsdUBLQ8nYmil9NFDFRS/WwYt8ETdP7V7EeYsm604+e0digT
uMk/7xT2vIBGfhIqzdcZj6u236bJ86Cb8ocn7EgBNN1NobFX7bh7BMAanKckiC0X5ARyOjgijdvE
I+fASuaSxkroWxvDzGCc5vuud5EviDd0zKWfdQn9ypEaebC7hPVUOJLvmd9LrW74mDGkaK3U0OHO
/nOIO25UzcaYzwzQ9ahCtRvbJtvtRiLE3dR2oYri89hv5riY/wbW6IL0Vv8jQslQpr71gNrHhisD
4CEC7zTkYyncKFJhMMcENzA2PggvmVQO2Hf+W61mNIdhVioGVshIS/D7pOovOcQjtXRpGW3JjZVc
F9fPkPY3YY4D73FQQgshkkJeb/NGwtTc93GPyM6zvt9TJLR8Dgh5sktNoUUrVuxJel4sexNU0E/T
8vct4kDBr00z4HH0J3XMC0Qi3szgR3cLkJIQ/5wkO823BeeYR5tbq/isPquiB+YmdOI9k1E4O5OZ
Wj7b2d1bMxXquCeyTUYqmWfKA7vbZYWn0y0B1KfRgaXrJPcDvaXgalQWkVknTgCvPzcYatX3AbYg
8rQOBLDlhCzHTh8D13vkDWdQNZOdp3U3YCgnkU+LMqtayHh6u1J0SbbggaMtHu8yjmJBi5FQBihT
Xjp+vYBxY5n6gaiwkHAJEc9TVUcdjhiVCyaES/WD7xwFsfU61KarSVMGGhr9wenoANOftsmZUhej
I5pfBznTigru7biBB0Q7KtploEDSH6ycagbX/jT+dCVw1OWHtr1TShqy/wF8iqJBdMEU2tfOVFz0
g1PsUY6f1EEskj2KQlWrNYeR9hbopVh2TGiciRgn6ChPYaFdF92lP8xL/uHJiMgZzPRo/ef7a5L3
XPsDSLBoVblxAORULh+t/HDEeE4niw3TvLN0BRSRBn9sckegw17rH1CqjtbL1OvfDu/vb7mQn1Vr
IEDNxnyoNIfDbmDVgJ5UH81JotH5xoQJoVDJZE64AnTNUTWITsnm9NFYxNBvf26kgCz1b1Mits1t
KZ7sHAv41j6hklDhl0+ttUExeb0mbAp0tLfhexmdrLrJcAbV12FKL31bgTDXcxUD2dTiH3x84VCE
RwUMUva3OvdHMqVUtXEU68VeeceUDD7zfPwiaCWj4RI3veKkDMOCnMeBSNnvzQGcDDSFfto+C98d
tk3DGW9lhc5LKWshuAZ68sXMIAsq8nLIekpIF0CB4TN0YgCkq9FR21Y7PiRbizd/r91EYy22wrkM
K6Tx8uEupSdC8G24i0WTKrVQgaLZHFsSR4bVt3I6U1gXq56IoffuDsYDdWkKhNpKSN7TXrImkF+0
Rk2Bx7yPodJWc2jBFTsin/I/sZe9qF0aOBFDJdrE701TIQiSt+zybw3Cgu+1TVZOPFv0ubN4qzxk
3dQ66LvMXvAXfrmYrLosGN+0L0kNXd7+QbRG7jAltRBE0cd98gI1UZsz/WzYioradNelzjWDNq10
w1udtdaxIhXZ4AyoN8y919VYgYEgxgu/4GLRnmGsXbzBCT4S8SlpK4rnNVydaH8R3DMFbknkoDT5
sqSyw5ICq2vfhUmg84CRnroPpSpET4jerjE5Qfrjon4TOE6xxrOASu4Tz/4iJQuftZJ7WnpQuRHM
cIsQ8hzf9vDghPlsF+O2BNRBhlb53vsrYkEGJ6H29zvIoHmeRaPJ6jQcVZjbpXwHhTXRd8Rn3DWI
sTWy3wUj98sRAEFf070j8z57UTSf3wKRKPGvJqZ//jfh/M3UvCzcLAOzYkUhOvNnz9k1hfJd0yWx
pCHGjGQ/BhxkubTOu9GPcOp+1Fe40FhyPH4s70lPOB2srfEECJBVNSYDsT4XTHeaJrUYRSh539al
wTEFpfljKliUPQXBxYSb2kJhbTAKydugOcLs2HdX7/nFqZgcMFMvxwdYJL+7rkyldH9zQ97tSnvp
q6Mntk59c81D07nT4CQCzABdFjp17rowwXLPkd3+0b2nYTtgf2pR8z2LI2rqPE4EokwN1EikYy/U
3910lFJcc5j1VEwoBLz7wIdDHqnsUhzqpsK0gvf8IScbq6YNHCYmBTfJitAt9BMD9Pvqbq2B53yX
Yc9+Jd15efDJLvRkdmvwpLC+2S1tPssUZG6j/IsUq0DPsUireISk7O4n9u/Anp7q0MWkPKP6ZNLk
5d/w+Iaj4JfSm1bNYiFc2Xz0P8O+QuC++RPO+MIkPCDySbqiGhwUfyGq6sTiAGq42miFl9ichT3A
fkyp/FZaDvZxZDd6KPLN494Ct+ktsFhMI4+UmzSzkmmpam/gn5no6hLZir4fysOzDhkJiO02DRKX
ztv7MFbS1j605bZzKLP3z5B31vgCUQvyb92sjjTlHiIW+i2dh4wjq2YcuhTNXCr42LspQXVZjP27
x+uovEl53pvdfVioBYSfamNY4rMrmUC9GRIbrPHnND8aRHWCZK8GMNaaQGfBiIcMkQ7uAtSvTiyo
8FHQSP/6i6r0vQBdmpmtUO60zkL6YIUcnGGFjdZmTqCDdEJw+j8NQd8To8mbz9lmeD+K/73utFr9
l7J3OrtB76pcogeFz0V7PsV2WRzJTaVQgW2ySmOH4GFvxWmtDjGaZFB5a8pxoK9EqS1vIY2OeZaW
J1cqsdOadyKjDKk9vCQjPD5knxzofae1PembYPU3y26TC2zObOTLpw+RrigW3Kaa+11bqwXzgu+n
7hlkcWMOjLaG3LxxFmDg2wu1+iJfn2zN70e6Rq+Anx7a2hJO+3FovxpTyjirukwDHz72VpX62TDW
oGA81oJ9DjdK+M+2LofTX/EDL1VeW8EiX6lc2RgILMv8iglxsYWaVnHxcBxSy8FEti8lbX6A3+pa
Bsd4EXfKGu6TT/TJv32GrKvVk8HnCEVeV1/R8cgfRaYhqpnVVAfchtLFTHWduGMGOSJGMXmY/Z6O
Ed4QR3ifVY6KHvdhtoxcVxVS89kwT2JGI+UKs6Is2S80BxFXHPJB9dn2WL/9Vb0tkdmfPPT/VV4W
29cF8v3LnJ23VrbvNRxfRolj35FQ/YBu8A7MJDseWt8v48Ai+t368Dlx/40MlvEUXLMc8J4pHeP6
TfpcFxJqze+z1g2XM/JZc/u2BQbEkkjnYrfB41YVMf+JReH7a3B2HYKkKxAz4ihATnMUEVlSnbMl
tiGxLLLzmdoQy0iSjmaBWsS+EfhrS0Z66oKwEDO8j4rvNO1sc8H6F0Lq3SoXsOVUFf3280iXPL/4
SaQgyFLMWkAlNHixoxnx/3Z6XMGjDzyJmLoaXO5uDRoNfR8r1HIQnPP2TGX3Tx5+T++qTuXGQe/d
n1D9hNe2bzn6rln/7iK43sryl1BqTxwI1oohCkGzUnFeIBJUy+3ZgQHSdjzdDhiO5NUlCp+Nh+tt
z5dhYx2aY0vxppQ46y4qcHhl1XEkcrxuzBan3alBrjRkT82Go66r6ME7qM+XtWnlG6R11qgAiM1n
SHWMlL/LtQUyZGh/VlIjGjQR2aY2D6MbqAs+jbLPnCK/dpJS0wBE6mFD2j46PqDsD/GURlcfYNQb
eNEzHqaEp9icWtsUCUuwxK2hCjB7iQRqcN2u6bSJwjTaBy7g/xA23ur+ZpLn6od9o9qWUux/rIaL
iLS5zhJsIBCcp5rd2kVvrZMLdMekqVGpprpD5CzsY9+ngIAama951q39tz6vN3xfS2igGD+Yh9U8
hXamabaD89NHFwV76pqFDlewJdrGGBjO+dZsGQUTSKnyZO4GurMInMfmzrAWE/tYRDDDMIuDqbJs
KheCq6Ee3k9ChuqVMTX3GfRHKSaaoYB9JlQzkSUzTMbuVVV2PPsv2baXQ3xOBffdWvw2Kv7JBeju
tBX8Ah2v9cChBSJxvFXweFxxIh3Kr5yMVbOxUu1EmUX3CONY45tsYWzmSBhsbZR6UXwuhxC7n6Uw
cuSJy0iIYHPaaeMZSYifdLX0il9/+Dg6+UuxDPyp41Zgz8225Httj8PXXeHyO0Agz/Lmi9S0kdJ6
oJzMBRuRip1QZQixK5AEcnsbkFiVqegtV8dBp5HHOSy3wEz9jO4YVcBkhRgrhWEX9Bd6773t2kM5
jgZXKmsjp4FhZB37k8rsJIIiTe1g5xHE6pgDvExfbERD+NN/o/wjmv+b7AkRkrA7G7MGGXRerU7a
5JrxrOgygHsyFZQqGp/g1jNupUQvX0g9tAcYFYpM1mtuiaN6Ue5K0nEJK2k+aj2ILn2zZ2uk1+Oq
FtfZbuIqJaVi1+NFa9RPJ203eQAFr038iyIOuBBLFPKBgso0aNipfNtYaXwpK92zsF4jMzfzi3AO
46EP7juuVhKqPlAjBcQrFjKdaMPvZT2sbYpYTEGo1C0dyivwfanIpIniBBV8ZtmaKXQ16fqKfN9d
vW/ErZxFh1FOJe45w9/f5hpbVyfTwInKSi3H90ltMGr4/mC8WFGcq1cwV5MYvDfBvNXA43IsdUah
6bKnb9VSKzsOq73p88R/yTacJ3ScTm5+zarV4IIDnqYRuHdAPfJsBUIvR1/fzDfdGlKXYl1pLAqL
L6+Sj1RKykasZkIlEPVMpmwckamcPpdlzOSC/bjTTyofN6N0lTE1jmejEJjhWSWiGz5IIbupX627
yoH6eH0h67ys3qiU8WxAMkP0IMKDoYN+jAEHtaNFxnysmopeEgw7CB9pcAofzwOd0Rpw9luretNj
TN4Qg0fuwOhaNHtQ2lmQ1K1K07IVqYojQ44wUjFhqTOOJb39KitAqIdRtyAiHmwYyQQVtazb96CE
An85EHQht4JxxdkOBYKGgYeK2cYWg6BZ05tINW2FEZpr+bM+1iqZ2z6QtmLk2LwPh/r4FrYZPtPG
e66kT+qskgncIT6/W3JjQHs32aFsoOnU/R3iaMldI2nYqFzCwO/iIEwV3SBP3TnHtlWphS4HMH65
azyltxgLvMTHu2PfrtRVoDTaxM1IwmiOQ1hI2EEREf5DLvPGTsDLQWZ7PKqHPy8ImHo0prynCcS3
6chYcof6ZseRCXj2VTCIRWOeA7fcVjbrcU7z5jA+RxJe0R5aTb8x6THTsZNsq+AiEjwlL0UDPTsf
Qz+pZ5kac14Z8ixuwAqv641g+n4FwT9g/B8pK2omuV0bYFBsQWZpoQwAay8Cy1tullk9yAoGWDzb
NSmkj1N4lLXwiCkZf/FAI6m/ZPF9wLiMMCWQf9adl/ONb4a3A62Ga7PEyiKh5rrCFWVPZgLuWTlh
4bBQ2AZfBUPfjGKYFgrbhGWtBgfL1GQN5HIOrc6OjY444pcDfMY9g2Qlsdt/jQL63waSkHiLLb9M
4mBonrYx4WhsMmTQNDBSIv5PeXpqn92Q5FP8Hf8mgxX+s4FbzjkPOnRJSBn9mD985mu/ew9vF+j5
sduFQMyxns1SOdp/UDV6XLJJvmgp/qwPcbW1kp+IvY4L03GDsGxyweWmF1ujTX7HCDvjUFPYqLxL
WxiODRM8WFlbfhSScRh7op77mKlC6QplfHVzx2VKTU/DncuPwYYXyvjzWLSipoMfrV1BDdlgH1v9
33iQC1cC9SKulY4bJJA/y7Z9pyr0BEzf5xJ2mZNm0Bk2Gjc0YbNIwWuPiYF0orVKfKXhVOi+f+IU
PkhaDD8xYQcTc4yz+XtA+vzVE2XAbUR1drjtkE6NzwedrIVFNNGLsdeXG8FZQ74MhKGgoAXmrvCp
b51+SJx3Xw+A/lYH5jXbjLBVzMAD+jXT7X/8eLFTkjfEybKJeWEfbgC0Chc9niapJccLWD6Y+SQm
vY5nEz4ZAEqYW9dpTTi6JFO9/Qy5QezzPLHsj3cXh8R/6FOCHEyju4Uqpw2tvDH91gHfnGZ4iB8D
iAKRm3AHIR6Ai99/2Ddf+8KHsdYqhTW3ApgPRRxEsj9hw69+1AeB4ua7PgIatTGakKy736cLmc9V
T7FN3Zt6ii/epAyBKUQWFoQa2MwH12+iwbPC8IACeray1eAqMr/uz/xrWmi1BBwLeDiU+J9Fp5dR
QshklG8+Lnsc66ehN78oSrblkrTqCEWHtVTBlam1up2FC+ev8XT0nACHbO4JZwpIrl3IV8qXj6ll
wRomLMIdNekeH2mhtbS9I0FEIse4ukO5DC7NNjp0XpmuQXDpm/uUpYcfV67xN4+h5vifbj5jmNLp
LCd2ZHqDsUWNV61Auc48nNNLv+7Vw21fmGR2GdFKG8QXEABRcmsQK18Lwrjt3qAftqvsQIfSfYMk
NMSGZpXoQbe/SNjFH2bvObgZXuZ68PJeW2o3ITBQDkQ9by18QWXFO71j4RHFB6bers86lAapxeTG
J9ZEJmWu988NRhbLCVPOl0lRqwpBAsTz99iMwzSKMLathvhd+fPsPp8A5CH/lTuf6VUpBckl6rfe
3WfvcKFODLMzd5fGgx+y/lircAxC+YOyXjfPV5A2N/EVZ5Lv/POC4d3MiLNt/edYAiYE4rtzAPz9
AeBcvTTI9IWliuuL+hBssTP3B0NFDYjGMNUUT7VkWyPBtOcx/8HOUQRD8fmrZA2top4sA1EmJrXU
uq6jhmFtHeCv0K+lujNHUiK8C6N5huARRkMu0w7jJyivfOc7VKD8Ea1SDdmqHjnD4pSN1qA+zrXv
uhaUKdzH1kOaDBwGrp4nDwNkm5sANbNqV1YykpGme7ck7Jv92lHwXJqjvbH3jsBzWkGsPNodxBag
p0UBeSHVZ4QeZndc2TN7NUCERCcIHRNzLKsapuNzSOo0CZpxGCDhfAa1mNrQXvr3O5RMzKnXFqhG
PPFQpefFmGf0uNgO49DiiGaSLyLUp3hmQmNeu+idmn01TqUHg+vyH+ncQvjnNW5WNu98CVHhAkkF
dug3sahNWCvKx7Ln5/PRGfSdaCkA2mPX5C7hm0GTXWnV7TtS7lq9S6QjRPWOqpyxeZp20tJNQdAL
SmN6TKz2lNNs/lSebBj6+YaKRargv7WSNYjxX2eQgzfmWZiVoRb4LgqHBuV+niGt0EyC7COKqTMw
vqfYeWZ96eNa8QY2fN6GCCp2x6tGXLVIeI9kSaer/jlOHkCkajQAUowMrm7/Z02O+/xPo0VTmODy
LwkL2a091NMbWiZ9aLZ/JX9KQ+nk+1nTBGOqPClIntn2xjFOyrQQbVo8mQX2nhSbgOtwa0fxHZt/
4aKU7yxVF0oG1cBUOFYTbK04EGRvMJR0QiEtUa7OKtfksGnYVQNI5VdV5MfL8XSgtBRXWtydFEmA
2sqXjtzP4CkmpZoKRw575Bj7b8JTzEY9sx66/5zx04U0JnTd8wGIkdySfQEpohlp/PEXt5LNxM2L
sbzYLENs1aGfMLluK7aBpMbkEdMighrJIV6BTQGvRvuBFmzRWH69PvB6FSpeC0hNNnMPJXzxVplk
JmEt41VcoXqF+dyQrPRDDUGmJQvnxHKiq5wICSqqsqhEdqBgGTlr1BuCW/EUF7tMKvQQ0TSRLFOp
ODuN9LS1fChH45yWSmKjRKAs4gfcHCjxTikSo6aCXv94VBZnMnpYloJF+Fmbg7nB99Jddc9l88Aa
khbip9haDji0DssnjKm0VBj0JnFov1LScDhta2leNSidFipnhBLBARjv/T7Z5optDh631xnLMKK9
uQ3nLuDXhTpx/E5sAe/DvdAmtR+di4fMV9Pp+YlBpFOGXbMfKr383Cadu6jsTl9+kzG32OpYrtII
xUk9GuSu5uunIgvEF50P6SK8cawUoD2gulEhGDEbAIqSBKJ62tsCRlX6lC0S0z5jqnC3cH3QlPg4
alm0GJDLeUxlmVuzZOIWeb8J9PXtku4DxCrKbSal4HFM5bIJl2NUVSsQdTbSZq20se9gHQ4yqelt
InDBQCAidkHG/vHEI6miUkedMEmvnhgMUanlpjiQCIBNWWC3G7o4cx90wvs36FsQb43CIgReU0+8
5JYMtj+sFf0NNU/+4ucF0F2SMMWcy+0bgEkBevY36zyRt7Hc8f8jsIQEWckl+PeA9ztBU0iKkqSb
N+NlWaZlgvRYgu6Oon6rJvUX+110Hit96ZdkYNM5YCyY7nbH28rGNCU+BhAKP41rHqZ0hKa+11H4
PHD41OTIa7eNzkZdERUI7lU7gcWi4wq26alX7akL4471s7JGrBOTjLdpg6fdc/IrDyr1yZ4hkY71
47NURnBG57VWdaAWPqZoEpTk7G75LsxPrbzuvAS/FxBWx2/VhANlnDVpHcMsFsncditX3SYXC13V
fnS4NamifF6WcTLWraK8rRsVbRTBnB3PrAPtdhQGlXqXe/I9aXlqmcDG+cBu1Sorf9bEEms/al+x
jTowUHNKO0mlJIgzei6PJtnv3n90M5JFjP1sxnWWC2W+2edv7pgJpCpm8/bmZbY5Bq1lb5LcGvgQ
QSVqEVNU/5ar4ocRghYTRcnsIvBGlFa0Ez5ReerRQxohX3ne9UekkfLjs6nz6DrNowZVAk3cK4jM
xdq6V1nkHtcai3lPgRBSBiIy5/n+YFxcsj2qTMoHzx6lihl3vSgoP9rqa5j/+VB35SNDeLycrHmJ
aVg/ZOi1y3I9gl9oWVUKmX7jubvtfwXLw5VOFVxmCdjEzuKnLsKkw3RPuGoQg6FxKK3MXqoswuFR
QHh7qDrfTobJOXAfplRo5zDdKYG982lBc1IWUKkogoBgrEoYVKSsB/Vn9a5sedNGQJReAYXTC37B
XkzrlaoyJAAYMdr5GUiGYtvuJuNPaRurNgj2P7FnApXFYd7orRcfQlcDhIQ7Ax2OWVfHf8jqrqmi
TVhNS9GRsiHcN3+Ti3HAj6RZuWkup9z+wm689RylBCu3KvO8dphi6h9FpIaFB+lyZ6JY3nao66Bt
9saawXAk4wRRdbVL5paT02pS5wU6CzW2FQsFmO4Qp++sR0BDYnIm5WusJXRUGvdGE/Lnr511FfdS
P3erasxm3iIhxb+g0qDtTFuYyH0lnXcXV2iNujPfWqkpF7ewF8NZ26MSLMIM5fS0kGQIGVba7cRL
EVWrQssbWq0EnvuFTRm+zQN2hz+IJI5TlDJA9qpBprJ9nrBq7XFtH23rfseeB/9yER7XfAitGUIc
kAaV/XLCMeUoIsg/FVbFjhcyS4YURzqm+3tTwUuEx4Ggp36GGN/zyMod9LOUQUBKFhAgSsWwcjhm
6FMh9Gjc22kvh4rivJofRvWd6Eh2Gghph517LUaXpTHuocOX/s55c8fYDmEsbiCKukovQ74J3QJE
TAIHXsx9azi8wcIlead5x3r/acAxae6URL/tSEFxfUUQ0r/hoMIjs4ZeiMQTklfSGNrd35KjjNpn
VA1O2qbs8S2V/qqRUzOzP81Np6kVCk+LE400A+BdGYoXm7n+4e0KzTakjZFDenjR3Vwlu/F2RVLw
q6HRxJdfVEUe2bxOJz8GmwV/DSONfHJ6+TRUxntomRQGP+o+jeYHyLa3nbQykgkdatshQwkSvlJu
jYPEOjd+hcXakMwwowmWi5asa3yB7OfvXVyQjdgbU53yPl+b65pBn5a4hkGE5cqbku2vB8d6r1Bg
gnFUreS9n9+kuqn4T8STugId7q8TU4cAr3Y2PX+HN0+bfVC6vlVcAKuXfPhOVID7HS28o8/7zloB
cc8Actg8hod4sZ1VpqcAQzbZ8Jeywcl3eq0JwOFXqrGcV1Mdhi546O5g//2GGuF61nljcsjb/Cr0
YTsNIjwv2Szkxh52eFCKpWnWYWscltoKDEkQo+1MrpD9S1qb9+DHvbA7sgSEg7DnPpuH20cR2Uc3
NE8SI3n+/SDxx6IlT3uQQ1km/2GXQbUlbwuPzosF0wDBTYEU2yX+OL0A/Slgpl3N1M/7t7l0V4YE
GYe3IpIqzHWPqTS6mSY9xTOO3f3hERbhZ56mTnJkw0sw9rE3ZO7ML/UE1c9ygijCBCYTY4dq84Uu
aLHBbJt9mJU3hhsJA58vgSNuX8802gpVpqs8tyBHcZvsAA5ij9bp63Zw2iNB5UZ74/L/MHkUTmha
Tna6BZ9R8ashueXczF90SjVYwixrNU9Vp2TWHkNhC6CvqvgekOE+FhJxw0vhnvTCjp8twNZaBhjy
sa7eQOXk9XplckiySaHtLhQB0ErRX8HrZi3hhya5LILqKI58narbfrLXkyZN47rnXkcKeX8Rxwo4
4uJkDfQ/eTciFVorwFcwYWnXPG8fRxvnvOu67LAGE/54IPOOnUyV78ETBKQDhBt2RPJ+fJBcjh9A
1oE8v6xlPAdFHsJz8v7PWfO1Ml64Mcw4XqQNFomXK3eBUSPaH7QvqxnaZv281tNUSVqXw98bMktA
x48G/AixAsIVqdlpcgxPeeVRH3jbVS9CV9oCguz58ktzuHDlWTqa6VgQIfS66dsaPg30s2AAzucD
yGgfvhis0F4pVf02EKQU2whgcnwOtXBiqDcYs4TZWwX104b3TV97JoD2MaKZPzqEeME8J8UwzPGF
IAz9yaHPNk2AKfR9RsVHRxCDvkuA+iO7H7yhk/S1uf/e94XymwAFdUbjA9mqg0l5bN4bavoJ2T3c
qbr/vMgul522mBF9Ero6MZx+1iewnUBQNEJS85+z0gqv5jhOg4jI6Wo0QUJRUt+zfAS2+8YWMWou
1eFlNhQSLOyQP/cJLcUvTnrBMIaLGQztkSuNO9aKuCaJaFLpi/6jCTXOfODMC9BOM66VLFftWVpt
o1VSLu8pqWjTzUyIK4WLoPCHj7TzQjqJtIOCpLcihMjGdbGrKtKrj6wX2u7VS+n/cVSY9FCuU1FD
2TWwFcvaTHDB04sHXUrmU4jNMsnjQlO64wA55Oh6j8E9iSYQR75Vsk5uGBrvxM5nb0S6Qeq26g5z
HgRFKSMrKCadI4RYO7a2dcFaNDOItkcNU6GOvl3tk/gQJ7P4Zsi5Cjtccjg+5kh/e2Ye9okaCQfB
lSHsk+yfKIJUH+dK2KuGXYCc1RZWoeVqzphwYiJ8gdqQNWA2Hg8391l6buvOenqWeGYIEFI8+KXb
qMn3gF1ZHWA+qLXeSgsFDwW2/P9E2nF+r1YFCdIuOKRPG4RwxRWLZa6s+Daaistvg3psbhYAL8c0
AmoR9lAs4TWAQcjgCSrSCTjNKyhei744I5f7HUNd+v8GzhaBCR0JBfLyctJu6onlJnk+ue7R85ti
DlQdPoYUnAHLP1ePiC6yur9mWRL6D0jFW9+nRisd2UHCYM6DA41LYG2kfLsb3nfDLJR2Y2EM1VfC
R7+pnrz2F7g2uKoqQWb+4pN7n0zS41HF01BMrmUYNbTkcrWAa/vxq7+h+q7zmFAnZt5hyxsjM61B
eqt5TkaIuknkvW+dTChNAxOPKjcvwAqqqKmJPOFzocfVRlIyVopvr1tQWb8jyNl6YllkDDCZzoqj
HMd1pCS9jS4E+PmVSsUj2IX1npKY/+OceKWLCJ13K1tbjnAn2KoDISAYaLIDBAecq8H0H/py7iAP
nPxobUaBnfWHt0lczR7w6WxjmnNpAFbUoLdJ4arLHrjIj5+913/5TEqKTpBrB2bNNg76kFya9YcP
boLOoWa/HVa8cgRxAUZ2Jg1NzfPBcGC6V9yUGWmB0o1ndwIzIzWv7li0LuzZxhcLoZakB80HBxxv
JzBlZXHEYfZi6lm0Smjvco/agWAKw8aXAfNN6AE7AJSK/5ESACKbXvVSe6rxS1DivzzgtH98pOE3
4BJgNW1p6PrhYrRRlMzAANqepncG4QjtjejByKQH75AE2kPifmZ4CMpAnFe5Wa2f6u8hsP0Qlf5T
x/oXhWTmEgqwG8U7pCvZUEwSVvrAn1f+7CnUnBkIBAsX7onoAA7C2z+Jj8Pk273R+NY2QBUCcavZ
fxBPjqcuU1+t6lbgSMpw5AB2OFgBqh855hHkzajzahlnyowqWmme3B0QNv6zSJxjJQVt4wrifW/g
rk5bgEwoMKeVFVSN2BdEM0RhKi1bd4FoSDGoIl7fHBbSh5iggbTzzQGF0UIpmyATHakFWih4w9km
YxKqD4K2S71/DS3M8oT13zhudEGf0+nfmfw5ElBQJzMXcnmRKSQzLpUnLbpV9ryQVkX+vswdVJz2
jhm00p6NJCyD2fYmmXgYe5eI4NEqIaM9E2ukyTlhfE5nbRYf+ejdX3zJJYAhYGab2+PBPAjujts8
hhGqHxrM5tYFT/YVhJ6GhDdt0jj802FfYki65DyNQf9WjohhbiSjvgFxbHoyFZ4JKhm1iue/X281
09H5ebfANoDzcLR4ET9cBjDRGrKWTDUqcjW0PCGQMgyc6SSlWe/YEt4W4f0KFYNSyiW73nr4PzQY
ditqE9gyaVog/Ge9A/6/Cs497Gvd8vvTykPjZJiYgEhqUKtOHl7uj0lcobvDRRJelolSDWh8pcDo
XCaAbMoPkvKjzly1RQwrFMiR9HYSJFqxV2e5y83U0ybJ58cUysa523Ek67GSA1PC3JV2f7mdIPJ/
5FiKY9MVMZ/nf+sYoQP6hSifUfKAvxYNIpEfm43YbCT4ph5C/EldZkElvaRSVPFkxMpnTjRgsm4y
GwOOw5QcSbHNDAxzNn5kEO6MAlxF53eRbSwLUMuDckRElTOUu7VQshXuSB3ZRrGB4Qmk/XGDAuw6
GOQu3GSODNrbd+XA5EVs60M+ZlgnUAaY9DNGZnWQmx3R6C4Gs2XAvApio+U0KrooPviTFR9mSAB8
K+Qs+5bmppaon/326JJrTFepwfzG19ADjxoEtpRXXhd3xWfM1W0xpIj3lJSIy7UvtKuurHMdCuEp
A6Jr6hSVrBTXHO/dGvm1sDdzwcVpHUPxbd3pverEDKjw4+lI9NPS4LdhruvLDG5PCzDsktN3kp3m
Q+YPggxvQrb7jZRDEAwbEp2ABDSqptPX8HpTY1EHgh53Qtdf1klG2qGFZWIVnDZDVdB/FqFK++0X
jmbcWuPOQMJr+qFOLR+T1kZMuzgLrK3Qx/8dJWm8tjbho8ISOzXGB9j9yBVw5X5AgWgi4GeSC0BA
nqQRZWUDshJTszevhTx6dHKcgnA8jbh/OJSSIiNNDw6n9odo4DpYkDOVbxP1Ef9x/nEeaS8zMseY
Mvv36CK1KaYy++r+gO9EgGj4y+smbrPoiSLbjp55FvpOW68cHdcj6CgbaUfLGxx70yaDLvcoVm4D
DyN03pCakKVmvJTfOFDya+ycJLWiLRJ5T8Z8uIjzt80HbNTcqhd6qwnkhRFei0Bpa6l0HFj2if4L
vRgdVMaCIr4j0JxROHGBrFB5SLNxWxPdYwbqe1sshMIkg1Mjz2cyRTiOXqukN5c5JMWBm//4mYlX
ughGYrlZfUpgfzkW5phIKw49bzuRxrDgPEQgNVx8hAcEYRt/EFo/L/753p444W2fbUv1AEKjoyam
kp6qWXz2XRAG7OSZWAb8nBl3gf5rwmQImmocMMQwRojnYG5LQtTc1mdrVTfsVjnHZQwlU/xdAtos
VXWt8bCJtaPefi1e5+lk2K00xB5QqUDxX/UUQtEer3wkd/YUD7kKPczfD3LoXnl6Z6gB0pJo+KEg
pMPf1YNNDlSLqN+SO6/HccvAoLPf7SDoYpQjINRlwUZKWxtwtifadsnJh8QUWGX3rpuMTBBBA3IN
8T8q1KHIBJgIwTn22TqSX7fXCHE1ncaO9MlcOk70ucjqH60dPaR6oqCqdjpDXRsKG/UOA/QnVO84
F0HeTnzvJa0K9ROoh7IG/EVs26PGRYIGByT8thG5fS0NU/Ru/6GlmnG92iLtK6MEy4KwF/ghNKzO
cBIAHStqUN5dgsV3rt1d5K85t8Hv2M5pAxKAO1TmSW/ZAf6Hzdx7P7sPbpxwax2/q3fBhydIwVWD
ktya86IZeaAqZJywqQLoIAIyQDZidskBjjWS/xJivGFfpwu3Wn1WOLNl8ST3YIFxqJoLWWmxc4QK
/UU0ave6Lz2BzoIEwXc1FVRzFXU8mCiWrB5NUc+D19Wd7ObmoVj+Mbq0RuQ82GO9kjZIbhmkQlkR
T80KzXSSECWLnd8tLkmOA3bFIPqK5T1p/Awdxkjon/NKg6wTTCLb03La5AhNPC5G7NluVvyy8WvP
TtHKadz23Bz4socIjhvdfhXWmM6WYRtrevjN8lyjoKG1PYJtj4ixCZWGQk9QwFUSZIcyijoD8YrT
KpyY27lclWnl1Fzl6WxgLCDUC0iDtZKGa19H1B6zg7V5SHBiblYdVnPGZooCHH89u/79bhWLZ/dl
1DrJxtXFvDvmMttWLcwYN20+917pxBQbTbP5HH7mXEWre+630D2wCK/+0ZWbprbS1tOtVKN9tEp7
mZ9YsRFH2PEuj5Jk3Olm9PU6wJEdz6/l5iyxpSfeXfbeuVzrTRJUXP7qDRa8h6P0RF+sW1k9Nyo7
met0HVjVBHvmR6GkK2wlH+7RJhMrW/0wmemZ/x9GmysBkWvFk5Th90nmN11RLiYlHGQPXZQ15bow
MjfFZ/NvqlYX0rUqCK7FciLaGhI4oqPHTbkMydsk3dLE1Abf3u37i8H8ZkaKT8dQACgqOeSQMHgr
tLxsxcFEyRPId0JNmhB30eD7kyn7JJzTgA86oWvZ09bNRrXCkYIlzJBZagdYndHPygN5YY/T96+S
PlnpGU0Yl9eZJNZdTUrcnktbx0M1wSqKdR2NJ3CuSD8cv1UcBHOgW8GAI6PK2svaXdWEnAc1rr7c
a1fegEyupI5yP5BA77uTF4vxEw9PjKt8QpHyt2WYkhesXaWTdgWJVgQC2lLYJxydPtBPDDxYeftV
fsDThmc1XrzZOxxbXiPnLqC1aoFk/2a8i2p0Z7HkU1Co8RqZaYNzj2t0JR2UNPOUYcaeFtEO3CAF
D/1ePVtbUxp+82lIiDRhvphwSf1YRhvYbYwLGx+17p6cJbvF/+1z7QTj9bg30zLx9VOOv2j+kXr0
6REHIDX3dXLkzpT0dklUDPthZ3SOkba+Gi50JA4GNwoL3+m5ZfJPsbU6Kc5/J8FLPlnTlTYbz2Di
AyUohtnyWZQl61fJJYljaELMc7RgPAkWgbpLF4fJEMTq+l+aX7KlXUj7LpuRwheIPzjtOUnsQXD8
BJKNWKA7KQaGZbLltCWUvvqVlDWX/S40Ox7Lj2TqF44aArvWHH6zrCnftovgp7wj71QxtHvRPE8G
ivGueV27Qde5hWwwsvy7qtYyNRNzuYhzVBRqsDxB4WJ0S+xupQKkJQN6R4v9dUU80KuFWYcjXpjt
6ZHKvSf2CAUheB1zZaSPN1VQxslX33PvPe9jUwAUfTI5hDbrRfOQZ+WMVkPLKmh9Jv+wUirMrxw0
OHOoAoFuMdfrUqvMkBRSLAqyq7Xb6Xh9/KiEU7Wg0tMtz7gxuxdNAb+Q7GEaw2eCrtTg3sB6+JtY
xLYnopizujSoBl2V95u1ZdARaIKSoUgO32gb6WOedFV4ngUjhRFdkVW5uiwmMoDquUkHQuOwZtSt
rQf4GQ/j4N7eLs7eOCenrC7Y7XsnNcyQx8ylDbj2kQQ4HpNdkNpQC9vmdpmQZbf2iEI77Q0b/W5R
Mb2XJ7njTPT+vCSwJbyc+Du3u8J5/lJsi0NilmDid3g3zn9coWoUfUZ1hH+dZkMX4Vaf8n/fEoWU
gyHz7xtF5z1m4vueJauraLV7hWbHBfV6BWu/9po6o0hGK9Et0ZLnMYB3kisiAbwHW7QyFw3OPXKA
6mD0qa2hhzHnXbQiAvTBEtC82dmJ+22yImcT6AWBaLnEGm6jzrjsOHt/HK9pFfclnvEY6DTWQPWV
E7jjM71A5nt7Gt0I1TeJVcGN2Iub/bwLfJ6jNCbmV/szUZCDEMiH0d+P8/QO6JhGei39p0WUQ7Jk
Rk+pRBP6ARIAItQuzZG+n3K3od4FX2D03Mr1WAY1SVO3JvGgiX9p53O6yPF9z3knnc3nwZ1KhljW
7pb3vbPT0kSjD//Kzqi1qjhH0CJWh60jM0lmZeR+C/d4meSjx2joE1/xaNURdZA2U0K0bYbDcgXQ
1cBluSkixldjkdP4gml0BHoysZS716aptT9K8Gl7x8THheD3f2+8+7EvQ44inqfdmNqssrHL7WZh
9HpVqpHYGmCNwm+YVfiFQEnCCALhHtyslmeySGcQhGOq/E64QS9H0H7N7v/Qr5g58060jahoAqjE
jZkZrUL/keHCqEm3GkeQNBWLL4plFkHfxxKbkrr6HtwOUkXKFobwWewcuqi3NgRjGCDGMKOHIBdP
T34oipfy0OInn3L5KAf/czf7BsnJegQlyqC3sweKmGJmpxVG9yZX6NwA/IG1TQK5BRBvzLfdAgJu
LActS7Nacsr04ZpQZbhQKBA+26X5gbWJ1qPdJbNVl5y8+TZMKRidfZaUaoe/fyyrISArl0Vcyf6+
boce52gK03XXRiQ4KA14pl8qMUHdzvdx/IOjhXNMbk4Z1iBP80z/Buo39h8AaIQWU1u8fLk6tNgk
nPQFlpzL0bTyzXVdJHjMg1n+DqICVZn1nL5aQBPMDNN8qYpw4Z7PlW1FS32wESRLLYpQCmMK5oKW
LwGxMDrNjz45fOf7KcNLbFyxCr+XZ/2m4+v3qxha7b+OAZnbZY9Wb105y2B9NQJy/5lP31sYA3bX
NtBbh3zQczQf5XOVgmaJATISjpC8Qhq2B/b+YFR7fM7+FhpDR0vsAcsegOauQsDWHTzZzKKXHtHU
Ah/1UEvnSBexoI5wsOnnlT2+7RP7orzoW7OcpISJBu0G93lsxyVXjsNsoNcalndO5qwSgTdlab7Q
Tj4e3T5TSaUdTjwfUh8oI0qp+fn5X33J3JGh1OGuHesI2SU+aHGsUHRtBoAOhFKQBwJN4l1bkyZy
fKfPgA/BD0+QmLA9tabaJIipcycGjt8BF+96EBlbIXTgNMOvXlMOOO2RRwCQiOcLIi0zTZAwmQuw
G38yZ3jjgFg4bVuQHLCUQLyJu+EyGeRJw1QE8eLX8Mx34GiaSJyxQYYaZJRC5gieSTRYYDJCSal/
9cIOoBTHf48AlOKYoysSDS3WhQW5DtuE++Ui9+0pKre/Z+kYLuZvDQ5cSMGR+D9PocrQumKVkAYo
4D1nhPX/tU6dcR6q/fcbFrD2UUnI2cnIFn1SD3WoVYK3RGjyKRtjxxbUPmRMoh85+PzfKJuzgV0m
cxF5Lhez31qu0g2ZeiNWcKAg7DNJBFPAqK/D2YN1qTitakOVh4/YfLdsD7fRl/IgIpGn7pVgbvmD
JtU8iVWS1Oqd8kJz1zMiwvTe7nfiAf9moaSaR8NMTvsnjsB/tCE249pPuffuBwfOoBl22MuS3U8c
JszpFjLdD4IlAXhdJ7GLX1K3amkvFZnB4VmQKDQvnyAWXJCVKN8OznYeZ6lSYAroAmQDvfJCQ/U+
kw6pRbkjkzTa0oBxxu13RUjDCxvOKqsXCiXzrojXYQJHf6SPhjVc/vSF+N84owBOmjEfWL8WpYU1
P0h1n2aAkkXbhZAf4rzlYC1cpH2kiA2NDw6N++KxcLewyJYC/baPr66g4a6B5nB0APzEtiQgeMir
kC1j1+nKPwkhwlIwHPzJWBII5cjtSR8FuzJShxwP6M6yNME/AxSyI1KZJN1YCNJ34AAatApqhjoV
6rEGK+ceomqEpmMmFQMgYvzrM36Do8SEsVPSv1werAUOXb2/R+S9vG+Vzwi3ViKFltO+zrIkQKwZ
eOQAzaeB4ojocL/AvzChSaJZFNS+Q7n1g2B04rj2jtLwow603Um0hC3/Dh+bN73wBy42JobqEIa/
x0dRiW2YwlkYf+MUzNb3pWMwVpD2PceJ8irwVSBNDv1Imf/tWHuoh+CEcqbKqHhIxg6fZjv5DxVq
18ZHaaC+yG0TLI/DXctPbldVh/eGHtahFQdxDOFVQmjW8AUGqEvxmX0uJzGxpiSb21SHumUlkpCZ
QHRtYHduryBhAKq2vEInEVPL/C91NdXS9+qydjHjpu2Rb9zbaD+MM7iga/4xF+ZpjJwdA9XCs/10
TivwGkCPa7/6joaWg5oFSr9pijNGwRdUzk4YnRthLJA2v/cEy+QfVDFjSwfTPZHb+eJnM0U6GtOs
r452iU5x1UcKntp0XIQtWf1MK0Jf1RpLby8SSAiIkm7uNLahTGz3FFH8oI6L62mXQ47p05MYTFIO
aldWscQu/Yw5UKcUKjWR8oBle6k5uoai2/pQWcs2YgFHvuxbJ7ATBkabgZfXkigyhxCf8f3jUGoM
FDUV0QjKryRXUajx5OfYi0szLAZrtaJVmm0Qzbfl7tecSp5YiTcD9b8fDKEajrP3LoQVb7QDBbIN
IbXFnr0z9B1REDkKcOhgm4pOMgk7GVtjV/thpp4P+RpBYeh62p2XAPxqIzeWidSTTm1ZL1/7fRGW
D4NEJ0vfJQdX0ENKsflqc0QoUEvemjIjRv+N3Rd7csJvQEzR0ToZKNPrSV2//lryYiXNJt/xVMYP
GZTEpuadfG8Ua/xDrMLEd9u8b5J9EhDZGAOfj0OQECP1d7nIijBRvOA8qKFZwGgNfQz49iOtQ60V
9iOref9K9pfVwbHnOCnqMRdc1JDPTkynt5xST6ImCRl51f928v7TSANXTUl6L3qDKPDomfGuHxfI
cUtgKU5xdSd6UgK8taPJ3EISQh85brt2QMQORTtabbqhxxV4PBRJiEckBUHJBVLXgeRd/GNfMoEs
xdkgolRHIzMqrT+Qg+TlXRGl8L5SofZxFO9Q5OiBChhKps4hic7u2zmR+Lov0XxMUj690aP5ZeJ0
qAiQrPSEJJ/f954HyWCpgiKjLC509Olc77vtOa/mWz5zyrkiHekKNHFfH10deBeodXKg2bkCA8Z8
CS+pS3CzgOB7DIfok3Uk4LPeHDrVSTeJfe/+UWYpDgIFHvUqEBxqeSRXgA+BREt/XP0fR2sDIQTl
FsTZXWTONyEdnsN5Cfi2n+FVMCO8MD5zPZbHx85B21MaOyiO48lS92YQsv5xypyvhLD3IgoaXyJd
ggEZO9DEiGeehO3ru7pRKvW4l1xknllKcfusRy5LSQ8jpMREzytJqZgnjqQo88enx9bp7hh3QTXw
JkonHsOUZmBBaLdyfT7JqKl0nE+is0igUfimBtFBRgtmBvwwyw2hs3ME59TWok7j4DriOoBU+RxE
M36ForZwyQ71pkB08er8Az/yKV6jHD7owLnmhChkglAPrA/gKaDGR83TleJ/eURIjRju6Z8j2fxm
omdBHwRueSVJZ5Xxm4jLSqJXPDWOh6oXDaa4W09OJaSwNnFd/BZ0bkEcLVh+33bDER5qCbjD84vN
5eveDJeqfdKhw1p0kXq2HFxiExTflegPh6bhnZtdeIOXyauh81QeEDcR41VeZH+FGU1fuf5NcOrW
yo+FjWaUmln7LNmGz75zxzFvvx3fEdKegBrHw/eV7UGmxo2Tu8AOkynDbhT/L5chU/i4Y8Q6hTkX
eHYHWgtL8m8HvLxFeooOOFlCbr2vpBLbJDjLhTgKhojiUcHoupZa5Oxfs+mTHwSESxcmOljzesf5
LYYwhUzC5pPn5bUzRO9R9Wh5nkRP2CxhNObLboDuEN4gDoY61U3cL35CJ8KYwFssaPqv2AOyJBs2
XtRCDuekMG+KuRgY23hpaImReWyoNiOrEsT71D1VVrjbY4UB01vlH9m0WXchfTfJD+pJ+zNemCpM
O+kZ7o8jNdelDA9DU4voQjED4BUvB84fkmtbp3c5iX5pC2FR4X5bfTLWOK3aEj/bcj2PwvDBb0BD
+3i/N4O560ZF9ECx9e10x9gXy6Yy0IfI61o6ibUvieCkG2unbUSe1iwbQaI4zJp7Bsn754M//9Oa
AyCxANIK7ildchql2hts5I0QYaj3Rfy+F+KRG9Zo/ZYo/oK6ntHXwnRJBc0DfjO2YwAT39OJJfA8
nAAsg08lCDmsD55wxKdRSq2b84p/t8qTyXGfIzoGOh1rinqwvx9xQLfUIvaYjMSEKbeFMVlYJ1lw
30p2Mcok8uefGltpb1yiobNvNtsU7MvftBtMD91aG8dJmL5fYJXaUp5GoUEIoUFbiBSfwBb0hTXx
uZmIarc0H17Suu2UYrtuXGIr5yicUNRNEguT9bPkOeejIMQgATqtSzQS2ITVG8VqQXjdFELcg9GP
pNJeBDwialBE4klyM9BB43U+fZxoIZ1312za58LHd2rBCHmuTv4M6OTrERJze1IfiOJdNO6cLGQR
vOgvrpGCtUKsWaR+3y8t9dn9aNidfInVUsrx/8IbuAsAdHk6dA8lUJ1otBfxfYwcIOblvdGduwFK
rexh8rrqWhsy2YJykFkNZIwXI7xyUHcD3DRENL6Iiw5IAh+1DG01Dlsi0AUam4TAbJvw0tKIRjEp
ksXy7TYguEW4Y80xI3Z+jehQVxuP4lKJd6MehAURRt3nuNfPeRYw/OBryZgOYxkqZ9eKWD4gKSHm
+muKclkBXwQC4n1FFDhf93MAUtHn8NdLvkvUrTIEqx4WygZ9DS/1flAImhF2uzR8y9cP6p8kAFs+
SP2m+P9uP+LL+1j5fVKc94ydGWI/WFNLK+oyZw4nafGS2Wa+JylDQ03uKusqF1Q0PvgZ6PQPH+eA
D+VtqnTotPnc4Z+UsCu/ZP0/NLwRHSmE4/0O+oqdvnDazRMRCuaeW2kFP4YMHyU60to0u+JczKKI
wA4gViQydnMlGfBxU2Am4vh+45mDXydRfYsJyh2g+mBBTZHRB0dUlMhKRx2TtBOyvfU9O1kTMM5+
BSYdo0tZnxlDG9AsOsXBijDgUHIO0LbiWfEAOg+Tz3rQUaAqEzqTAfj0uqrO2VnVGmo8lmOJdckJ
FMYK23It7iQPEvkTBYZMFNgRYQ4U/2z9hNYJAcklD35DKR++KpCBCcMVdRhtReMmc8oInsGMzVtc
3xSS7Y/2gUNHWYoNHZqtkQSojcnH9vWNek2BRYobJYGGGnqv7lSDPaedR8BYZyvhwzvPsBzubZcL
83IHM9Tg7wEQUNVjfv/y14ZUaKjXvIOFOliWy3xa0opXR0SVYjf99To/6suIRtnAYXqsXn/LAXKS
IgdZjBsc22qbt3VQNOr82oO5igtvgHkh1IX4qOal8z+iNEnWKr3Ydh0J/v5q2fBzfn4HTt0Ibiuw
AqUtrWCJF3XbwoB4/5wkSrwOQeHz/SWI2KzSp3fxwURXIK3va589oMPLHajrPs5m/Ga+JeYJc6BG
M9ZlwtiQJ54GT6TdxZsh8etf6pZD7MrAYYffgvXo69yrQJuEPpOC/SA2Hy365mRk+1C8j/voegqB
gJWvLp2pwlMwxF7xy0SByz6idq6AwAZRFzXP2b6RXiIpeyyxBlMVzo20w0Dr9wP5ggH4xwuDVv4S
WFz36+QNTTbgjhXt0Jx4a2gqlBPXyx7y8JZIIsP1QbTVBsNavSMh5JdJvsrST7LmK7Rd0YHEaDte
v3WgoaDM6Djwq0IaRhrIA1P8RrHj8n3wzLqpwZHJ9d7EdQ+C9wyyvQergntU3oPgOXRo/18kMJMn
BlhfZ5mLqRD7IHEW73R68rdc9d3kUVUqBdHAo1aDCYsQ9TLZq8Up4kArLys9a9oPYJYpInVPacgE
5HHcTKc+P//ItqjoB4sEi7srMsrR0ghvSt83zONdS6rXTpK9/T1TKBH5XQAOu9o9wvYC7ibs82d0
oxZCME3LcEEv8T0L/j7CiA3QhDmj8p5HWfR8RV/W5pZn9mxQfCS9geFstdbmamDHN5Wbr5ui+ZCl
CAqhonHcDcT9lZ+9dor9C05/w1+4meMi+nfeAhb23ZWprIEjoxydE3f6fsrdsF/1Z9+DsGjUSFm6
Sx6bo35AwyJRqmjLelZ2KiBB0f7t6ivf3mwSbNWQlVdVogDD+93ogetqqLme66LvzI2sEFiXRIa0
T1pG5/mRWvUlz5ASDhSGl9Iz3O8//OeVZ54jG6BQbtn/rwphVcLcp9gdqR/fCefYjpl6MBrfkZJp
x+NM0x264HREHhA8YNM+CXyOddBRIz1dZayfH8C5pXJDgP8gJVS0yw3MbUwoKQU+5yeypkJal1iX
d1cIs/ceRP3k+Tq+8vG/K7WsVjc+5gLzDYWk5JHYJvlobXjQYVHbbR7ltMuDxRjWs0/hwmzCXv8/
GBVRg5ylT/LEujtRNk3xqVdvJTbSIDeszq7aimyFEM4heYkV35gLAU8TC0l2HZXFXwVC/qNdj9ZG
qxIBj3XhPu3597iQvC7ucAD32rsO4cwtsM9nUeHad10rAx1xs6eS0m3zKiuNW7alTwEoDm3K42kx
3u9JiCzRq2eqw+tbOJrVFw35fZSqyCricFgA8HkHKWeC3xXKEwWYVWm4rCsl7FK9Sifizmb0zCmD
AzhJKUNpHMWcRR0esuMKzGd8fTY8H62JLaJjhNO86jJ+aBWTqSeGNfzpCFKVPlH6oYegkXBkdZtF
e38jOFs7veAkeUBHa3T+06wGCsKygCGjs/2H+cTE/nK/ON3gaTilnwKF2PUmM3pEoKRouc/JlPy+
oiW3upnEVMnBLimMe/Oak//huKMfFGYvh9jwvsP6y06ZMteEODvXZIPTLc4im6HPn4fUXDOntkfV
NV1RaLAH6S0rVzYC7YRsJOH4W+s8JTWRz012bBVteINUGTVJl9TwEzawIFOIoTSF/5DpdaWuy7X8
+jABd21fke4/OMwQPDBuItJIhERJctalaGfD7eKm6BE8yuTn7XNsRVx1zExlTPOw2TadIH3TMk4U
T02dl6ursKWT+avdg2XSVZvszO1USCnUBdME8rXcSUIrsWMnmj+APIgrd5kQ0Z+jw6kNqohNvPOS
5oKhqRgk5ttfV/xy4wgBoQgGqgsOAaiTV/srmtaoGEqx34kNXAiNtX0cH7o9TJqNjtGe0rHYAbVH
KkPVt5BQFj1XXBvp6qaI7PuNCs2pqak2T/NTUKhyiVjF/MxOy22mR4ADZvcTDKmkPSa19ZvZJH+I
ct7tG8lpMSNoKKgXf1dO5EgxWfxxiIDyMEDkxAm3nN1CNwKPDu+Z+T7GiEivSETRpyjs29W96XuH
aA7cUHDwmook4Ta0lsD3driLBz3tTLpBZKf6D+k5A5MxTXQbzLOtt2hEmSLcUTwu7Yw2iftY7Yc/
2EtlYi6YfAV/KCkvyDLZjwiX/9xdzDrD7KDkeFP6c/quHFt5qIjQxkOVefMxugp34WtZ6M1ArdEn
/ETB9j2G2o4q+1xdloLry6Foh+kJcjbZEPLqJnQb7qiPfs7NUXDvk/6JtWdzWSDrltwpzGrvALMp
VomJbx8B6i2X4SwJP26ArCGKlZ3EqTscjS1JiZI2M/BF8IlaiISrjenk7QixFngAZlQLTLE9LCEP
dbMgsGZQ3dEeH945Ez4840cqMyZOZL4DHn/TxwWK+NL4jNDjxZzbLXAc9jflXJdBuBdy5+oiAW0F
qY2zxisZ/xCXRwhUsVr+Ib+OlOsZoeSxy0wVYgwbT9Jt5TX/TR2OeGF5T2E9QpdIEMHJVmrWqCVK
YnJo1TmHqpyggW34dbhDxcMOCh9fS4UrLqWc2s2ArmMZGAWaGO/geUy1f9BtaZZPmevaY58H5X6D
qGI5e9VhCL6NRHINACWc4B8XguQpsYsK46ttaiYYz3Gb644EsKq8Ew7r+BavCN91QqF1twzHxXXr
caKQ/h4aSMOKkG9bNmYxRzkY0j3R5+GWdRjOgc6CM58FWjMNWgSOEnvhSWXq9G21cJBEA9D4hY6K
MFs9STJs3W9CQ2Yy7/ecOUtUCjsoatUxFNL/EYvFl1DByCstAHPqB721pn1OyCsWqWUtp/VIrhfI
vv0G6m5pzW9W7rhJgdgSALc766sO0xrWoRfr773K7s0e03K82yVR8MjdU6Qe3Dw1NgTb0X7u59Y7
idHSJ1Q1sGHRo7+bsrB9r0s36d+h5VCU/ysXN4xnTM2xSMptecXhqFiVSEyY7mhACL6Yv4jNlUhW
MTiTCXi1oWLUYVSuLJ1lN8OFVA7P9ppMLc7l3vLiyE7XNTxNwxMHJfvuXzmz2BB4kmECTXofV+zl
qwazdH8Ak0A+5SomOJFAn7HK6YgSRur/JanfL1BIJ6m1uQWV/5iWCTivmvwyB2FXZ/vSjffk6kDR
X/tsxheck8zORtBbgjjZD6vFMG1H2c9XSZs5NruP6fOIe7VUtxz8X4E81BG/hIJSAj1v36W0qiz8
2mrAPRpX6xf2ALCr7Fo6Bi972vgCEG2mxaQAqLeRGk6X4VWO7dRoBpzMFaQXICs7aAq+qBsjlUJk
TTnPAxzUiaTJrroW9cHvNsLE8j0P2q4ULCH3qCIJhMrrL2dwin3nTOBtOznzCNQiq/iqa20s7TDJ
HmPmu4nuVBlO7EJJl8aT393B0jlQyNlRbWUJrQpqTyVVUblX7VpnabGd69p7b8Zw9K1Ydp4SxIFG
/Lw+xBnKLZwy9+1+rI/Hoz6UoNU444tI8NbVAInCyome0hwi/6/QNBBRWtgLrHvQSKIOfXo3EJLX
r8rLik1Xaepd9G6Cvp3CDQGKVw9RQiO/Wv8geDqxAxnsVzwzcpHnj+Uc4dAHN9iUf5oxri94nSLa
YE88BXuyDrm6MdTf2ueZqvVe+o98kB/9+zc7i/9sP+IUVbQ1Sq3DYTAgC3IO70jlJWR3JQnKa3Kr
X6q9rcjci9Cz/GN/NZBzh4qtvffzUdS0tQ+VZ+pY6wKO/Jwa6UZfBmXcKV+jGrUPDCsRs7DnuPRc
GdB748BQ0iBVFueJDel5Qh1SXnIgE3G1kTsmVVv9t7jAqiuxhVSarVndp57DJJH+kZZKYoPMFbdT
bFwNH4hcjlC8BQyI6lpK1dR+9p8Y90L5bj70vgnS6mosZnT6S9gQ0OD6g03ZunFYE8c27F33c9Kl
SF5EVfwz1TX/Zv22xIqWHaGDRe3wjQrm9t948O2nQ+9KhDSwemngkebD2emuh/uKBUVSm8QqYUKf
IskfGuVq4X+Wkp5IuI7o4lSvN0m0CfQbfMRK2dF/iBkjZXi1qvC2X8WFAeqDJFV4CS7ZwmhiV/Et
AFnWb7GXmNzPlWbWsy9VUm54n70W8rCldq2Fmbunonue0d9EQvbQf3j4feyPOODZo9zmdxDM9V7C
vFvGRc5yy5fQXFwVZrU6lkkkqxmvzaNgFdG6mawP6Eu16ISlDMhT/dFKZMKy3N1eJ1N9S1XUJEb4
2pESi35bTSk94FmgfJ2OiMC0mNm3LEEkMKYXCznN+p2u0f2liV+nSreICHw7RSFCTc71YSRTcnrR
KwPzhajDKNlSKKCwsXkofugz7K9zH6TrTmjpTpiuZVon9A0undpeez7wJ8rDv88y69mBdvY+9h/e
yIZD/HIqoZeao91ihMNP9xo+Kf1KXQrnhsGk2Ev3dlhA3zFJRS0HTqDut2rEGxdsYg3AwLqkK3Do
HhB2cNoUZ+fXFS2pRoMjnj5OFlT4EsdndJhGt0OBpfCxZy0B4Bln11dn5mayOSAwdCY273u7Kago
6KfskYb8/kw+wF6y92J7UwcvIIY2EtMWOQlEmfvxxRk6reaRMprPm01NRbAvDxbGVk8SQr49cVKI
rGVUAk2zupeCY/NxZC1M1ev++eK9FRGu03DtJw23HCd2pfszwb2pP9ZZcl/Q78WLLKPxh5psUzCZ
qNQeC8TGTjMjeMHSUHuOIy3xLcmCp7hTUBfVqzjE8HDXxtIoKZsQhu9bl3OmGnKG88S+EtgMzDl7
yoYMqOvOOPN4RNfZy26tyWF3Su2NIECmn9NmCNhK0dv0rfdRWyLDtV3qkyeaP5N7Pp78lIez3Nh2
cO6ZSiUEcZc9/HTu2CWoreTi7y2skfD7UdASQKOkYdhLw+mXQVX1sr9Qhlq89RUUVSlTyMWmRvxP
E/HoY7+Q6pDgsYQHX2U3re9bg+AEnLNyhNm+EMTHCf13SfHE5k85eWeIcbn+zgq0A3yyL27s0U/2
j4fsRs8Fxxy0NbhAGo/Vyw5AMhrkOsqOgvunQ9B4vddnM1EbVSvOsFJt6VZa4rVc3GhuvBumryBT
bSYdiUBR7I8OKJra/iYgZF4USFCsMnptt9XJrVezSPnbaeobt8Lv6mucVH6dn74mROu35SEKtaue
f06hvGS4FBNIoEVJZ0LAuD6B2LFWbPrmL7frhec/cGw0HJX4NI8u1Q0rYN/sZrHnB31skrUSf4N2
WiBcz/7OLifmA5NpVrXM0bJXKw4+yt1crASFu8h3ZJ382t2WfXaWM1jx5ATiKZ2vRF0XSNTeGle2
8EWlybBeQ57BCy89ysBjcpns3dm+oCXTaxY7UDBpyOj5q2tNSaEztceOqh1Ywc0n7ZEzxOoLQkZ3
KorFb7RUdaYRkHiUHO7pcTitAlnrQInfSB8zAIIHnRS6EUKhUg/vhEXiPowEX57FqE+B9H8KlhH9
UvL9JW7/tGr2T2hl2qLrMMPyVTxMW4/6bIzrSgy9Wwo0PTxsd6drEeFCpC3PMBveqa+YNpdYvJ7C
0ePDdOHmFn/75nxgo8opn5A93H3+EMcbZWc8uRjINCIvlH0i1P8QLH9aFlRDDVKKjlxRvljyawqx
k9yT5KEWRS1r7pxLX8eQLWHGqu2kYfkZLD494nvAvGZUgskNFAkEbpwHWGv3A7FR2NuOP2rEVbdc
Vm6wCpXtIlwRjbUaosNqPz1InQ56Cye4oXZ2AZ1uoaW3ocMCLAL8XSWeDDuqRPUaOlj2Y0GCXKao
g2y0KMWybTjbLB70xSC0DZJwlyyDhv/o6efHZOGbQ17TlhU5aWEDFMCAhUrNm7kp2cM6Ka3ZQTst
hm42vUXLhzx/L4RMDYJQTHrm62cw2Ndk5xdMMlywWXg8df5Xm516KA91816tYmgFfJBAJvr3WdMC
iwGWmxXSThK9WvMgbqEoBrRmXa4h1vuMVAkUV075gpbpv+5JqyD4Pbd4NLwLytATtUqwHi4BI84O
uD/p8pxfjUb8ZWJMcQk3s8NmJc04q7LGOwpeiaJazVtL9Sansw0j4td8c6yXom3tB6eJJQySw5MR
Z/jP5dZbITrr7AUDtNWhMoQJ4caOyrggoYcK3sL8tmBwiJsl+dZn5WaJBYteuZbv8WC2xVdjIRvX
fVVdcUhLAwaIf5iGSW4ry/EkYBw0ayRS7BJx/+9y5rkoLNbrPFFICIoq5seyvBtAkZi/+qpA+Drc
fP11JtrwcVqiVjA0aNRscNiQzKr7q1tig+b1dacdFQ/T1RvsanZmqY4AZx4RXnqSvdfh+r4wPWjQ
KpwokEdBsH7sLFZKxiiYAutUlUT8uorz+XlYfsJvcMXKOFrXbKN1PplJEcug5QleXg2aT6dZb0zi
dMVTqpt6+rTt4Nl8dKtV9a5evY9+QHcFzuK0jKj798r7SHtWYumYmmsAe2uyBYU5JTiNdon8fbyb
A3zecr9bOo3NKMASgYw3OZI/WreoLKfNjEygiV0UKtOhPUB+skutTVySUOycFDj/dGYgATRDJMCY
8EjJnVIbFNK4zjjuyPHHVi6wjimgTBw2cyhjRSwfaXTzV70HEyBRqIekfmi9FrZMk5XaNP8CHh6H
nHaQ7QaMqNkyx40ChKGxmCTqneN4RYajQv164s00P8do2BJ7tYHfLGp4G7KqCif2LnxTyIlKvzqF
pQb3jshB2YghavG5RVeqLXnnTLSy7uOYKqsH/yq3zFlJHEoSf9KSd9w3GleKw7pgtsdTc87FMgyw
7n4BrjOUgQngGKGDinvjVlj/vwrYopTw74M/ktWPEQF/WFKfy5gt8F9/hBsmligHfdrEAA3p524V
bY+Qb1UMbijvA/chKVfbiuUDLNgP0ulFfV/FU+d+CZNHyFr97i6rHJM7I0C8lbAn4etmvWMr6SU0
+ay9N8Cd038xmZZGAZ26SoMin29WonQI+uY+1549meILQ5Wviw+OSPtln34SZxNE0ypVncNfxRJQ
WG1apAQLzuiWLdQSl6uBFaniDS53DNxEKgd59ZoTsmCcCyfwH3ySH4aLfPD9ZPrBDvzQ4VYImJri
G8PhrOW+pxkOjDkCZgIyvzzFMjX1Wsr+2lXGhwKyPxFBJ+VhFRJpLOSD63Er7Po+CQbRxSzk9aoM
vb77c7Fcq95T3096OshnFshFQZUhmL6qs97snkYszRxADNh9Atzxjf5L7W/v9Ew4f1kAHvaPtZ+t
kqpnCpEzSINVs6ValfDMQaAsHOifqw1Lv7EaEq9Hq0wtuFjHhC9zN0J9+FWaHjpM6rd3LSkC2mrS
6orXMPLgzvJYYFRoAAIyC2j+H65R0gYATeuFrCbEAjvxt4gFjFAaQu/qAoEqr0DBbsa/YVXzMG2I
b0V+rrfmZbmRIFN49VSppkPcxuWYcokw8lJ6glT1J+xx1jBvduSlCmDJb4nyUsUJ9ttbo7cXCvu3
xo7J2H7ovhY53JcHZpwGlm/+hyW/GdUBTOwDNC8uY1rOkuFAlMi1DsT0mngJnEYBTqsPLk552A++
3UqJ0INXlVUnJ2KC0Tcmm23HwK/ESC0eHPblgLY5nDhwKhttaYC1kyQkJ/OjPX3MA6gpK+4x0H9r
nOFVC0O6jofqYdtokl3SompzPqm4YVU8roaihdAZfdZpsSKfmtMkQ2KNuABxcVXpNo83qI5v3dGs
+7zN+RP0iT3h9ztFNXTsPZgqe4gfbizTMMuk/sC+yqiblKJafYtvG7tFO+KDTZ3FcrWVBJln9C/T
ocAjkXvfvVLZdeP3VNP0JclN0BQYQa2UCZVjF6ULq+XaHEautRd2Bprhn4neKN2x4IA8YHsfdR2D
9p2ND6JVY0sDz679t+hLGhE7fgr1RaVvdcsSRhaBWHN5ng7Q99chiWyGXjGoTiWHEhsGdiDGoPQj
ux91SDKfXc6W9D1dS0jnJvJ7FEnfS9Mau7lic2XUXIF85Tv/FDL+6vXAJRHa9ja5t9YgY/KAJDr3
ATPVI61My+KylaZH7JIyGXWT5u0G4oHTYsuy/9PLpjPH0YPxtOTk/MFG4GWoT5VyDxLrhu1FNgsU
sBLR8kPVXYAnmSeWt4wue993IDaCcoAzEh6+VLaDK+u8TGg7ZFxuqAy0ayVSftGMiUJhHvs50UrY
ey4wS4mfpSIiwFLd/kmZC7UMifcZFuhmBHdPvEcuQREWRXuSObDuZibl0mRwcfd/QXL3OHzziv0E
QRdeG5XIXKphs3woChbpVMEPpDyC+ilp09o4XtYbVQ3yGbfEOUsuRRbnbwlR2ye20D+GKlmitYAG
CUHwPY2HBG5IntY8cpMMshfza7LdQk/d3TJzDQwh75s/n7DBvGLWjLz9zCT/iGDySusidV1RlRih
fdrWccoMGkX76aDmalJNrn+sVhw1jlAkxexys7L/8+UVIDU1cE89/39PraKq2bl89t2JYpWY9BxJ
sBLB0GJtcgQSFUxwiotjWo9crvqFjr7SjfS7ItlWUDk2hlYMuPLAoFuV4Twe7jGueqe3xZJFsYIH
Z6gzs28cT8lKAycwS/9927Sg3Z50Td0Wk1M6eGMBYUDbmbYj4yfdM5Bt//Xzk0N9CSLCptJvgyFA
CJuO64OUwbrZJfj07UNSqdEhqYbyWGel5hpAYnr7/IprNQWqBST7TXBauwroXsXxZguD3Y07MhHc
V47+3DjLXT49hX4z3LVNYGP08QtddLzUL4LbK4pVIpfRmVSVgQUEUyuciMCTFEwwrp4MOGKx+z65
ItpxoomlUnmWP8rvwHMRgNMfb8Ul4Yu+FjYxoaN/Kgiz5xv2iPlUq4RkM38FifQuav3skuGUffkI
zLbrGJ4NTEjzfSEXCzk35r9SSmMRnZOqatBuUqHMkwdkHUOfYYYZdxqrHiA/yMyhRxsmLFyChYM8
puSLbQkgAsjmNhb3zsTPe+S5gQMlvakbkutJ734cRWpjW32phk+3c1sc+WiNNM6gyen7Ciy9cWNF
B+YzHSLWeEJRRin+wfFswZueeUQINZ60Ie+V5RdbXiOUSuQhz5LyO1jn4BdBdbRZix3vyN9PsHG/
PJWQ//ulG5SCEtNt00DdUx8vQ2XknIovwPXGVKZuqOdGXYfNRVTWj8UFQPdz/9Zws9tqNeiPe1dx
olY0aeLosdnaHd0xBEdyvWtKiEqIti7NSHzMTJamRG7xOTXlwLLrst4n/8WMO42EVaOJJPOyYdqS
TiwXqktivzkpX3fYYbF7TM2bgY//hBR4vdRstTHbUmT9CnOvUSu3t2KUmMOhq230gGY03dwmvfyS
du3dDstUm3QXFx+urCisLl8qnviBBGofLCtQ4J1m3rPkgG4F4Qa1rF2EoAR7pkLnTtp4o7sVGih7
sVf/yZ6t3MJtrR47JjyP0J+bqtiOLipYRGpVGa1pgbBir1kcd+4gamrFIpnaNr6m4xX0RcPRVwy3
Co2UJAS0yM2n4zviWCTTxtjLjCM5E/cRET0uMNFd/2/J5zefVB5hboETLdUnw1ylmefYvLyqAd7i
GI3AnWq0kTOM8djrU/Clbj3WzpDi2KfZpYaH3ERbUMLNyyZZgBWPWl1wGiMov/m8UbqPhrPkJX1p
63zsCbnkFqAkx0JecNP+yr6BMqrUGXRZaLiSeH7RXouu6gA4HeB0+7YDETs6uVFtdfUVoIZntuGs
ibvNmEm4U5+0dw2ruorYesCYMikBYCOzO5z5sPG3dmMPo2BkVcw1ixysa8OXmsGbkatUZ5C0FELa
WiwEfQgdyCFJGl5bRwz3PMIqEmS01EmZQeEXT3tWtFOAT7A0Ote8fZr8hJwwFgiLL4WsaUItlUHp
kYJpeKd1uqbUoxoTx1RHoy7t7mbobV+wAUW9Gkw7/ZMOJCq1zCkwH+4hHZzwRLlpctiXqHwSbgyr
ALSWHRMCeOvVvFUzrBeVBRhrhL15D9BVZFWvStdJFoA5AQCa4KH3v7DLdEmDFiQv5bOXQIWBFW21
8r7US5Jf5lDf7iZffWuiY37nBkd1fdipX8lXBZdzJJ3ilQokaz/UtFiVP74so6f4eOHuaE3UQMjJ
oHmq6EgLnq+wfnhxwBWhxxKrQxKDTxIme2/pEHegTLjEirzvtST99YiBULUNmrfWvq55fmz5ZnAH
wi++fffByGqfE64kJy0Q7myVR8WBoM+moSFnMO1EHB5goh8vd3N3yzAkv2HbJ/RIuN3DxhNbGGEp
g929oiO/dOda62aiSs83Ka+jh16eTa+LHaEAwP+fkGfmbnpdK8C/70kc6m96ueVp+ZVdi91PrVeO
uvXnOFuMUB1h3q8ll5WHWdcfdPUiPcxPPkjhsLGnCAl2NS+9vnckllRsQYMaMinLjMupvLVJ3AeD
u/vGDcImEb/lTCnGc45FrjQqaYHnZnCJXVPykEpEPPVtTlT6SalM+7LxGevtn2qB6RYmk0LW6ViB
HblhDsac/uLQrpEknMEEuu65xtaSPSQhCLLMWsLULo8rYqD6kiZCr5GXOf2wuRBpbmyBW+vN0UHO
DL9dVlfGjmx9kXTdri0GJxm+XfVkgcubeKO1kbMXRV95EmDbFfH96xO1m2DkKkuyHE+Pp/15hdCx
t2wscrR43xNiXivPVe5JaG7bjuYcT4wBI/A4lflZTj1Zq5D51FyJuvRaBy8jLb+KEHSLUZlUOWVk
Qs66nwlG04/Tovwefv3Vd+H9Db+cWNxfpoOiRlCmpvf09BL5kN5MTvQhZHve1DC0d5mq/1aRCmnY
FhZGIWkHbnznYQ/jEZl4EjrDSFG8SMUSjJNJtMkk6BfHlxIGQKZicJoi3EJEvxWuOrl0YIiDqxgN
bbrL4NJkXtaAMe6QIdQmu/XRuYsjTQqm2I0drc78ZDWpABZlO6c9yorEc5Tw7C3qLXSEJbgcl4AL
9C2Sy5euS1wPzXDqTjGIQCl3dMyNH+uGWKs4k4NH5L8KdvBVIJzcggdfQ1trWgxQNLT/pihK7dMW
qiQ+Hb+a85z7WLUx3MXWV9HYqH1CAoJkafpMuVygSYomgB8ucoU0IEaiRAt9Sj2KC1+Je3Tytgw9
safdZbAwmc+MeEY/XcSB8WlCUmAjuAyxi7Snq/g58l7rHrsoxF15rBl2vrKzhvPwtCaxV5SKvsSG
rJZp9WiFAQvw9+oP1QYuMgrNE//PtUsBjix6Ixbw4voZf7XQ2aEfRyPb2Ssh1oeCBu6rldWVT+U+
9MzX/MUu+/kbXFjdBtbUIZfID7M6mUM92NS9JE1ta0Z1sOTfaOrdqYceqizfLANeCyJHf/kNOrIC
yZ0/nGNrr5bRdzkhq7NS60a1GYEyHBhPFFSAS88xaVnT8GTeVBx+fZOkD6G4WL3tT5YMldtifXBE
BBQzgp29B8kU9sJ+xt0nM/yISb23l+pB70LjXLXIqGz1YBhl6VOlVSDwUtvwMsVMC3QGeNg2J0Ms
tGVshkjdTUj3aJbKRnrZTQ83zuD/u6XGyvUlrD2naYN/Juh4HZBP5H5f/XjTO5JsF6waQ0qnr4mP
XiSvfA96rdV35xEAu+agmU7KhMAFT3iI9c2zcnntMLFcCM1zXjygfEo59NMh29jCLsvQOTP8l6Io
/J+LLhmWYmPqxTqt7Wz+5w5VKq/0o6ttGA0EWUdsJfRYOQnJ7uph7972apKNE4EPtE38fFYId7Cr
Y6v8bLeJjhmOA9FZtDIeEISuezLnKyDPDQHq7VHcXhZygpNbtndHllgJjAONPgyrlGAicn/1KI63
80jHJXA4TajRGNvI0qJnvZIrWhIcL5PIuEs4Db06bqbzOQNHmX34QjL//VaCfduO+ryLuB8E/pha
2jo2ASub46EdbawP/NEUNViWGPAvdsaZVYG+kA6maSf0cphaLv9szkFn5vA77LY5Cc7EMHTdjKrY
Qzqlhv7EUikomBCKJIFylJLfagtnkOeO+DhIplTS/dLAtbWgQfaXzkz4M/W28HdmE+p/Rb88Fsas
lXA2qyqt33zrLV5T1XPxLQqJyu3ks90rT+RNSvSEo3JiS6YPBE+inXNdWrnfZOylPnxkbUy0nVfV
FPm+ZorwHRdpRu2vwwsFnGHBqzJZ+W+imHBukG1x4i2HXKEDswz6QuMBjBI2j0omGxFAXuWuhd9y
Cfp8PmWyDsC+SW18Bt0PDHOuB/gepuLleRxNWRkGi9fKyMlx2DmlkCSQJJ9AkxQIIjrhQgPuq4+Y
srWsIpsUg6u0SWezALUVizDH0kwChaZ3d/t7ryvRVD3fHzBt/dlkMUM7v0+KzxfRH98ysMFj1UFU
loA9A9IDr6y2hSRB/NYB7xLMGzI4bNv+xjfdy8wCAd3BG6WdZeQ8NqLzbKBKW9P7dGNOj6qD4gZz
swVRniYgNwsw+iKzkL1fnd6vAcq5wMMDtbgLMqVw3wLjYw9dzEFIstZgL2rhqRYmmKkl6w75TvF6
7M5v+R/PeOEWtr1nBdQ9NKF0XdT/Cf4C+4O2NzYJsQwmF65XeUn84cNg3L2sdGdY3y0KTbMUeG/j
ppJMsyqbqlzbEEgdLIO9OKt/ggJeVEW9Jo/09fQlQUBTUl5EZo/Xty27vKRSdVg3/578AdrxbSRg
ktsfcnXMiXCB9C7f9ZAB36eRP7HrneebRqe/LKFw80zIAMwFwLsoHNAUcFnEARIfeW3ADkePmDJU
0aZ7Bsk2eciO7RFG7qXN3F1CfdvkC1Cv6a/S8A5nc7ukMrqGoA2hTBMaW2yXZVzmZn4CLA3WC2+I
G3BfCxoOTX1VhR+l0e1fkZY0fBz16DvHQZ7u2WjmrJY0EpDYeKpWfQcFdId3Bt/um9oUOH8bWKH1
lMS3+8zrkVwoBda+kO6MIqCLpcxwEPi1z27V6W17MxlueQ4F2GiGg+bjzvWym+Fkj3mfRsDf2aLS
z1xdIo9Axb9q4zH9+9miwk/y/XB5qrTtL4jNVvxy66Uwf7QgS5Z3WLOssCU5wjIjrSU4o0rSPtk6
S154OXUVs1ZiwMBP+2iVtLSK4FdSU5i3GkMB0pPwDMYI13ruRzjoJLdJ6kSsgbMCuAMAKUbxkgV0
Z7lM2RDK7N8Vf0ykgDZQHHG7fmYTyaXAw1u4FGd38/6UUlzpPb7XVnj0JkmJS63MDNpFOGCm+9TC
EC+AeU2b2Y9faMnGqKZx2aGfWkEJqjgxJUvWqjinIEaxblma8njseAQK/dV7HjErntMLs41gFY0g
dJUMYKiS0bmNoUX9rM9KpJ83eEpd8gDRrK8BZjlnevAx0L0GVY3kw0UHzSGdsp5BO9IQd7A3BYvG
R4qzrQrwbZ/rkTBEPdCYBW8NaE6d4dHHaetW+IHQUW0yOTQQXP+EYeaQuUZyzMy8d38XNejJiip2
8MUn1MW0ZphuPSC++xyJGe78vFUiO7cxM9utFgs9qyti8MFY20Ed6rP6wxWuPvIJQbNhYldcb3L4
pW088E0/NQKT9k4PoBsYzw0vLN+jXqqD5py3y+BcjLtBBhaUcKGXc4kOdgYsZwS0UQKdOrsb3QJt
zSN4c8+8gFfpIuPMLDOvg+b4kkcyoIhTCdlTCC5PIetXbF88E74QBBO3G4DYZDelOK1/m2Wik32u
yfsh/EVYVUTEM9A6UFYB0SNmjnLWMVTKySD3FiD+gq2xyNDuS4RuMtsajeRYYfWldS4KYpz37+gK
CIj4AzEwDFnoBWzjilx5gMCZ8tAfi4DsKeSoK9m2ZL5gxGDkhGD+DhpSEQMQMYuXCCLSpslNl0hr
cmcWJ2Dmvcn2NBKbXPvQ8JdTD2YGVYRfmSHZLImrIWG+5f4vRmdEKokMsw4HgwhNICIjDkULUICl
0BRswhnuzOm5nATqmgiPZaxyI+YTKalYmajluJvMSoLGccvw7cIvTfQADZb6nQNRzMLZ9CdcUn/x
0mu9qFWfJDmqBnle6L+QQZha8pm2ynvFfpTCH8rmnOfs6T0NI4XuGZPvbd/QSIF1ids/KLNf73jF
dzfRO0WPl+iKyOr9z9h/Fy2kemRDINIpK20wYsE/6k7DnkKLhnuDBT5qFTFx/Z6zgBw3Jo+81gs2
p1i2dFpKfqyWqhawSm8RHWfZMIYKfimOwfMVFG1he6Z7FAE6uZom2Po1Xr3gzOneIxP8K+ZqQXx6
fKwCVNS6Ozg5cf33ysCCuNlqr2rV4QVOHcmW4A5FuOQj0BFsTGJAmzlQKQmR2mdEOJyH2xKXBR6C
59XVurHH6C7PY2lUdFkZuSrE4lWdIFZNgHKH5FO3+si9QiQjwvcFcbvx0L8sDnuSZyYcUUC0vIZt
fH2NkZEtBB8G9ENeMap7jD3sFXYD+j43sTytpxnzbdyxxWcQVDnfcQjV5DklVCstJ862i72qiPJe
VxuFNmfEjycJHImaYpYC1mcl5I2WSwOXuQb5uX+8mHJt2u4l7FxR9lOpJ9EB+qoul2IMt3pptCp6
tzge4Wu31FA8V3z4FTPzbM4Z9cor5cpTgAevcFv6l4E9lbcSXDNLDtLa1dI3qs3HAjquItfrBk7/
ElG9EG5zzsX03ZBLrHjYBUVQFKsuhnkgZwPfKS+Ai3Nnbwbqr6QI2BfxOXWhjNIlLSDOohoqFHmq
NGxbdxB9EptI/x8t8CinOu8q7RJOAzJps7OW53ZTFmLzwsXHzckqGCEPwBUupVu0PBpfUhiAqRs6
YAbgzN+FFaTOvMlmcCskxZR/EJfZxTcPhEcjalFEg+9fTpesp0aERWhnnd7ht5MNLffPVYfs9B+b
VCk5sHBOSxn5Bq9A/P7/ECDaabg7Ht113fMK5SPiS9faGRo5FNd5fRVAsMLoZ371Mhzh0uy5H13g
94k5kZGFopGMy3dXKOr8n/zrl/iGA44OH9q/qMb95C0DlV6BnrYWwB8AaBzbsjiTLgcJoPdaqOw3
/uJflDUPvQ3SG7zeqg9iuF941VVLpK0gfZOMNq5xlWVeTWlaN02eFBHXHb+mCoym8UlOHVqXoX1p
Vx1RtwfZRWyor1jH7BA/TTheoG5W2Pm/dJVhLUiMAmVkzB4FJyQXmhGRk617M25fj31O43ZTutxE
it/8PXMnPd+W0x2n3bd2d6WJOkY/9ajTla5SIAZQ70MnIc57R1aPZ/HuJQyFOLZSEuihHg9D8EGG
7TxMuKz+blcq6eYuN2MFLsubTexnFmSxKKRaBEP/QswaSZYTvzBYMAXlj9aWMrdU9CzIUmzVjRSa
l8UdIXUsQLwgU+cRvNKT0Ex0NKzjBmuvWPXcTYWTR+5laq5oRNpedx5wpAkniDdcAgfWx3A+IalL
3ZdefBv8u7aeGmbxytY+pTtodvT86guVKy6UoO4E+Z2cvkcIlSh12NkfQKlrbCktzboSHZIQOQ9y
6Q8b372H+Fx7px7Y7MQEshv4prv4kFW43Sz0+ivQsoGok8R8vDwsj0UESfZP1w8tgNyma9FjZFFf
eVyx3JpZvvPr52mKWG3Zj9ew6tepbhLiLr24qmjfaykwH5kdYVSqwlwgv/nXmWNS+26jw/8W5TPo
1ju2seI3UOJhJGa9wHlvolCy3CEQgJfwEYxl7QgkHcFwMbhrpso6XqLbivY6FjUOoEzampDnQSK1
HLK2ah/ovVCj+k0sRXD06AtJXh/DIPFlpXSJBHMNIWH5s57LRhxfu6puzOFKsB3J6ZXXVOIM4ZcG
kHykdr361Mtvqkk2ETwAGaFrlzJPiTaxL64zUil+qOpDDkPXtIpLEmiogAArA5IwtRbGpAHC1IbH
nGo296+U+xcswpxh+ZwabXbIDqyW3X4NBg0ZT27Xnoma4FxpoNxZaNuPBVeT5hU8yDl/M/WO3I4R
fULYhPIzAHKIunNnC0tNjRzMJ6NgrTp0GV1Y+qIQ9miMDUX4NaNP5FcORwxOw12r36SeQlqsMPRG
pJNcdC5oCbUGko5A9jtyeq3nLK1MqngmLMDP7bi3a8HWfSWQIrvcUviFGE4ZH4Z5Z0jwLQUqwx+8
LXr36+3+CV94ldl2HVZKSNB3BfwG+uv4Edn6Z8Lqp/TbLiU8+Yi58jt4sp1pQH1ElP+lA8apuEhp
Gyrhe+NEVMUav7gjVtyMH4vnICqEpcZqSlzrQ6XoclOyH2JgqhUnXFpApUR0CiyA71atD95L/PSs
gypeQ0gYxs6hchuJi7hIDFLBWvRkegGzab1vU9n0Su6/vypPt/Eyxxglo9WiirDj7zdNpA/mZCka
Gj64FQDp9KYDpz0XWT5H4n3M7kK0XO8RAkS2SqNTi1JJeeWSC9CwuZa09r6HsEZ5aM271pBIYxlt
grsXtb++C3rZkYEPJamzSh+zfHxHTt0gfyZpaMxrVgjG3fg5ds40ij05qrWSafSERfPrvgWa/s5m
gADk2SJIqe9CXjar9VV+DGxBpqyyQvXllzeICArC7c4DqVXNqVI9PT6UL0vTZxp9Wm4GyYHrB8GK
FcESLpglbs6cDxGKYHfItaZ0A86XvjRfN5koD6mGn0E6waDt7SFSlveISY1FH6O0aKBH5naL7la8
JlwJVcS+J6dikLrmEpP89uHdv5NjpekMyFV+fnMiJZs76mF6pnpNbdk6Ryv/lBOURZ+5jljUdelJ
sx+g9/UNl3L1lW7BQ8BU/QsWa+tz1RdLhAOLNYdM4EMuQ6ZPYF95YqNPOOaRm1f7a4y9F7d42f1P
/yTrU0HdTiUeiSpG1j99WW9j+RYc4JoB07FS2oMOuO4DD2Rj2Iy03GfGRfOSzxC4da0Una7q8Tbi
XOezbeqtIHI2yNaU1JC/+eLvI9NtYQUeQ4l7UINkL92mHj2UeVxqbog0d+sD2IpGZUKYs8v67p6U
FCcdwppHW7eIRO2zM1m0xv5PGB+fiiL9CYQhyv4ek6/HkOeFJrhqxbnAr4PhK/dnSKeZeTbUt6kE
qg0KDYIjq8vB7ChZyVXVi+LgOhHQBPzY50hupo7rJEaVBhdwmBXzcNy6UxIFfHy8HTzcmCt7vk/G
AnDgt2COlzWz0JxYiOx71Gb+M4kgG8m9EHtPkcYxtgskKMmZSYwH0FAlOdenEhFzqh64wSrl3QHU
wTGKMJUPHfCevGyrxKX4dml6U4gZRMYaxtarunXZtxqa4nYoAY5ERx3iVtrTOty47tzg3cqy+qQf
eDB41ljRAHoPw+XNhOax4Pv3/OSrdgAiyD2FTRH6zTCleCSWYXPuK0NMkErTqepeY+EAOCckjRIU
jqTloe7sQHU4y5VpokfFT3Ye9JLhP3LVwrhki5Pn9yXyl2R5sQkcIfJEC6/f9mPYqfKKj3Jkha1e
ysg31VnCz1TfS320xWAuCfloEESlE3E1EP5LByiTTRcNb78Hzmadn12qVsNe9t89gicFnVQm9t9F
wMae2+twLTNuSLInxF+lYkUl21B2X6UI7Xvarv9wUZ+uXYbEX6ddEfziYclhYM6JqyqgD4+bfE+g
kdb73Nvbg961mUvU9iF6wv8orK8XzMUzsHmnqnUxjoL+h31Y1rR3eND2m6W76ZRZx1j6J1t/7WDt
n5iDHlJjCYoK05bDjPIKKt1Iai7wcqRUTNpvdygTyjWWPng0XhwJBzYeNTr4fgN1FC4XjNuCNuz0
L1lVcVnqxXCrbaxBpaeSLCTYLwSTB3ewUAQESpuNaXxq6tVjisJE0UdB/fKqgvH7lnxySTlU3j1x
mnMK8iEUlgfzvW0pq44TjLdR/0G+FEkDtVICnCQaNG++XTC77tZgq8Gyuo185iHcXmPQRmfM6v7m
kbCqua01Fhm2+OyAiM2ICHVdJLaDfy/LPg6coqOin2JYauW03q6cyCTNuJKIznB/0rcCwbCytuC0
VlkYAc6w7ObrKmnnTztfPsov1NY4uxjfXHgJmg3ggU+gTYWMuQupcCU9Uyx2+Yqqywo8lou9hlEf
o0AxEZ8QYXbqDKaq1TmsUeucD5c5qByYwhiu4LdTw+k/xqG4bfu5qA5ns4FYpqccrTQv6YrYX1EU
2HCo3l1wdhQv9ldyiy+LI7/xwjGLExlMOWOwpi8zFsasvDVfbiqjpUhlhbp+p6iFAGVcKSgCZUXZ
UbUq8tFG5Cw9QqN1pxiQHAoAnmYoZ8T06kG/+3lCQXCq+R3l3CmZhCMF83JDqOiOlj1cCFF8QZs2
YuKcW8LeIxc3ft2Vx6D0E8laylzSkDscMbCUCOmgyjBKxniGLc9lRVn+UMg78VYe7ps6eoy03r74
b1WkP88Lp3cOX5bl0VRlbUoqv0xXlexpTkMPDpDdOWe7ThIIGNKgcGm9g5OYNqmDfPcsUYA2+qG5
JlHXGFJiOfydWxSqAN9YzIh1p6II1xPC1MXUR64Hw+hU7FaJwRD1VgMuP6l6gezDwMKKJrcZOiSo
d2qqepaEz1fv3KvpmtEStsx+NImfpnbBdkjETgjKGMjltf3zzh6rYCDg1KHQOnbmM19pQQN1HPaR
RObMSquxBoBBvO7r+KaI4i1Q71HA/D3MLrXANeBln091eA8S1GnKam+g04CC8nQarNOiS5vA5dMf
O73IXYFP2vodLEBYb26A8KhLq+juvLElIya3QZBW1SBOuvn5130kBETttMueRNYaLLR6BYBIQhRP
lBnHeHiJV4rMZ5QEZ+ba6r6JyXIWv5k6JJT36/S1sx87rdSxAZSj9XdKLgPu4SWwjUUk9GqLSL/E
VvGl8HXYgWS9X9NL1M+RDNredsHTFDZo+zpkXXyB5UXUGLoBfFlMA3CA+XjEn5qYQFIbQWUk+J5w
AR0KQ8WB7rywFH+Dnzr8rrGqyln9D02vGmJk7zE0hkg6kLFv8b6eqsb10yIkYTjNQ8Va45cCJRv3
UjtcbE4KiztuvP3V0oKlxi6HRrSF26jhjpcn2qylXxREZGCOMT2twkKf3C9vydIhu9ffSblfZLIE
h4kRkReGGJs50NVYoN96U1QDijqRAQJ2UQ3x04j0/e2G7b8FJfnskETiAZFoRIPsNP3JURtrkVUU
597f99RzkKJ3xSpKxZrmubsBMtLAXu755AVWFyTScckTsWhGfumwr+bdLbJNL57dTNrVIk/wehUn
g9kQQ6NrBmZoQlJumw4K7OGm1mL2WucF6G+GKhV4dsS60Wle1URJdlUf6DJowpT2cAQvEqIdSttX
M73ipLVvJXbfexLRaaIHFUOugn7/WAaRf+4yaX9MPpwsfVUAxKTYDsRME5NFb6PcXMlmmhfy+NzY
bCxXpbD4L/3ea1jO/muFu4gqtaTUK3awpRuiI6KDGTCHZUOPZdgCzAmtrLFYvmNePOjkUZ9uzt/Z
Vh3BhVNK/O2oLuTi7Z/SH+ShwR63ZoKA6yuX0FVQbkhh4hT0WBq4kB9TAOptjInLHbPD+acGUb45
y90b9zC20YHUp9U1kS+PQHoNLFHG0k5s58Oa+uPy8ZChIopvvDom7naISqVUb4hQ9ByvfEoRUP/d
Z6RWW2u5jFWJ4w1v5kdplj7FITAzecpWUZNBiUp0rqLIW5oK1B5x8N3/MWl0/4ee3m24dJMgG/5p
hjm0k2NKfg8sd0bcvgwgmdvSw7Qpi/cPp/oDopYUc4y5+YH+GP+Z4JziWGMHDfpxBiwd1uF9DO4E
Iv+hLwZFZ0G1u9UORFxRwG6TkUUy4Hmn35qpAqcH4s2r2Vc5WAFl2u1djm07ljOLiFibzyiAL1eI
uRsEyE8HrrkQ5EzOSDv07/agHxubbdh9yVqLL23GKFZzQp6c8VBZreKdom1n8DjkIA5Kp9Lvm500
swyYctOzLMnUlr9eH8HM2ZYY4kCtpTf1ruaCnsEi81nztStgkXaNbjNNQ0V5zvBYdTfOuKixvQqV
4pr1j+zJViAKS07uoxSa/eKhK9QRTBc9GBwDXaEuX/6nEkAjTLwlxOTGzeP9KPSIbZWj9IG/bbMJ
p4+806y2CbTTdOZVVEqlO8EWYBFKZEDYEBV9zcPRHksIt3TUTtf+9hryzjZHW56xlCl7vDpzWeUX
u/jZt8kR4mZQwCbmEUF4adoVQCqo3SdWVgx6ruoWKe6ykn6Bg8irsT7zBRXZTJWAEU5lZe79Z//J
OvAPnAEYZ83BQpvS+5ewH0+iDhtrdUKqU53hRx8P7ihDxk1g9HQWUSl/vUQ72crLuX0j41fJ+6dE
/cFuIrWEY+28Q5y8FIt2htWo2yEnkOshXDxcYWUkLEBZjeiCcb0SYuVLHnVKQqPGHuUe802ADO1H
pTRbgAS3ywm2AvA323dhc3xXPZ+UjCV69WtCVTi7nyCbZRbNneqpkZ1j1b8K4e6H5CEZ2y3+lFuA
5+FTyEDEniG63FKz+Rf1NODzoqk6NaUXU3cfQbgtQDfZDpkLTG3mCc7hdDiLT84OAOay0F1QGjiw
1SklOoodAhcx4RwKA/17JXJgnf5s6BDyIHi9O+hAAlI58Z0iX7Wvr4oVJnwoHbZFGEW6I5nt7OyL
EopqPSc8igZZXno9bW5pcx6CNGB/B9W5zsyg3b8KkoMOqWtyT/cLN67uVKvtRvEMR3d8feoA2g3d
dThNMe0XF9UQjnMIZ0R0jE6s/tcMvhBIGjCDY1CeOLZgKzfRKvOjiiFLqybTfPQ+L8Kjmhn0f2dm
t50FiCrcOk/RU4Wzo9QE06qqoD41DNWlEThxpAkJKb6uzBmnV3vVusnCi/KRLN6Qf9lp5YFq65K3
P/ZCBCq8XsBRpd10qHoryoK59AW1t+m1HkzD8BrRDibv6llVd1Kl8QjAmL9uhTN4FkWPHhTxNJu1
3iXMFgxOxRcJzzawTzUHtwK/7Usua7MNfWN3DmyRW3nCaePbN0vSOnkdHWgIbdwfs0dA8qqW0BAZ
ZQJKUG99gKfuFBnOVdQ2alj9nB2FhKLzGUcV8i17EI/ga0QnKy453BUgw2xs5a9QBLZN3oguEkb+
wjxmwnnF+0EcUctS/fayOA5MYs6ZbM/nIpLWjA2lfO0wBjGi64dsWZBl0tTBJ3fADd3psbeF4Xam
wFY7+Ibbx3IxjpBj8DM3G9BRf5UhYUCSKbFkEivpuOGZHMHtGxD5rSGKdEszrlEaogPrCwWBJwfd
C5QNWnubbt1jCZl6S2mblsjmC7YyFOS7OeC74Jxu8uhqRywe5Gtph9sSRY+W8Ek5DiV5UEof9t0m
eJqAMlcb3K1Dk67wTWQsO2o3PGDj5OltUlaaiO4Ba6TR8UoCie0sWpTF/A8yexaB6IY24jNSJcTL
AxL8o9LTi55Tw/ZzCsG3zU4PQGwE7LvuvypxEF51hErV8h08ES3nuZrtVpdh/qoF2dnv8xGK8OOw
aja97yMG8FZQWw8muX7NumM4FNNsnQGNijpZdxB1uPyWUHmZePOcjqoE84fr9u2fB5OJVrWFnp5F
44TYe44QBmOdj5h4SVUvIj/Zl/axPxrdS+RmEDa0owp7fB1XcrUtxV8n3A8b9K52hwpwlezmTCWO
95JgvpVYGW1/AIXP0xF7s9XPoi7xRqJ0yi7S2WjA3zemnQyO/2MtMyu9PPDq9FRaS2NAg4602pcz
PpyuZjQ+9HnzohMpSTeYGDAgvTbm9Avy6vV1L1GeezYzwLMftiDDabc+VnmIhEci9yNHyuHnIqra
RQ5ibbb/ZyUZA44IXQuwShkzZO2YGOvnEykps5bXFb0f8cts8I6jtRCMY+ljzf6lODmWpxXELltM
KSICg08RTnKcmF03WigqyRfaV/4P8fSHbrP9vbnYVHTPTGTpddLWxEPe15Xj1Gt5mO+pMl/lsN7u
QnIaCTFuwrPIRiknqtyIjBF9jJQA0NyILBXD07m8vp/wEJ5y8AbuJ9SolStn3xPYhwbOOenxvxJ7
DrF+9NkWcB8V/lSEMetC+nLUs8n7lGrQf3K+qeatz428CyBUxPz+1mi+PSDuKEbnIuBQ5FcszyKV
0NmwZbPjtJjreT913P+t9qPetpxNvqYLez54VKtwKgni0LQSV1laVFbsFtnP01jCuldNW2F15OgY
ULfluNFE6W7QG7eB4UdjQk/R4zBSQ/QK8KLqBrDgqnlfvFXOT6P9WnhjOspvDWsD5F267aEi2cST
tZSX5Esb795Is3vJDwRhb19Z8V78oYjyplswvq0XiZd1p3lsCHVXhvnz3s9ASgLw6nl8L6hasW7n
VfbA2o93TE+3/Kg6C1fOEV75t439mAmyDkbPfChFd/Kxn74ZllZy4clsKVxJumeaYUEvzbuKBjMo
F/9Aex9p/LwsjA+RuFXbRz8HVQ4Usk+YVF5GZlOufoK/XYAIG7/h861S65HRek0/mTvNUYwWXbjt
W1qZnKVftzOfIht9HVQAecsA0eD+ymCS8d7m77CDoHbNNCdu35+JEzfZ9BSjVbgt2vPYOHH3Dmgs
C+r7OcFs+jTSTp632H0YDvBKUF3JVfoAkP0mgGgUAphOpIgH5hjaIJhdHJIn+KC6SZSAyHBjdHtL
3rq6X+iyLOcTjlrZGQFEG5lsE9o1rIcZJwkkxjGSWpvkDe9ZmdyEqGgoQ6/WDrv0s6wrWEKODNYd
USCcMUnfweEnaQiX4inXv2pW6VChA0VLxIpz5UrUv5bCGBmNfFVEn8derDL+sjD/L3If6WNwHS0r
RKNQISTaUXNdYybDBdLyab2S1wwv0T7tJxWlGkpzS8daReNmnwqRBaFJ0WU7VcPqJwAtf1PcF6wX
ywYahS2B8IIfNYwqxcv7Q49E9Sa5qeuosDGPVMVnc2aSiR+FlJb4nZHhr3FerwR1K3pkzipEyJQ1
SISPwe4Oo+Q90vSfegyRWt0iAROAz10urXEBUKSNbMkvv5/3H4JRkdPLFdvMfMBSRM4CbYWYR++G
LnvRh9E8NBNDlBwBcOCH4b3aEdczBs3ToPS3cV81hQjDgw5uJxXwBwT17Lc342h7tFf/Z+G3SpvO
oNRx9noNFnUQzyf4AZBNMlX9KlPt6yrREYr675YpOZFkC19cvDWUElfATjE9ztsd4ZnfgvWsDKZ6
LJfzBr+CuKu4vgMa7EZngVbxS4stcLv3XxDUwe+l/1Zg6darpD3VdjGPz5wOUQB0brZB/i2VigAc
SwezJ8mBc5V2OPoF233mthrxtY3KgK3HfkqnB6yiULiF5lMzcC2Jpcq/COekPzwYV1tE2f9eH8/C
fglvsWap6r/HTU/sRJyofYWpB7/g7UpWCpLyAKtV4VJWw1GDzVWAyIqiW8/3KMx0K94NEIKtPOHl
57YEGc0wbso9RYL4H5+u5smkWjH++sfdlmMNa39+jbShJNJArKUrGtcVhBDljnoM2D6bROM4vRG4
5enWZJ0r9yogO6AWZ3DSgIc8apOukWZ1xoJRUEI1/XOa5i7BjlJXCCD1qvj4VFjZD5igQZe5VJdx
fggZnnW9yzFsOVbrM3OEmJcGtoao4rnHZaBuQHreLA4xJ+aIgMo6POVf0sgFY8TQJh2hjvlNi6iS
DfO1VuuqOUSZyJQtMWju+HixFjj5FbRfc+yKphK744MJyD8HPkx/6vMv4yIWh0ga1sS2EOsCAIs6
rlcoOVIw6ByVDk93FNs2sFQbv000EhPFAG7I2athNbqi/dWUccJbf7FKrNTDUXg6Agk5SNeDvdvM
SfCfwY6yFYOcyzmGbnEiscrqhCWE27vqOHS77PDIjA8LKrF/yMg4n9WsoNMJIiJQLo2MCyKVIjv1
fwd2xRQYjH0+QtFrxDhFm9FNqmCCwhfaJYvpE2fuFhgkwGcAEgLiJqoS160sPzJqEOSwoFmMVzEJ
pSYQ1DUOjIyV363ubETjAhn2d+x3DAp1GDnCJk+PmazhVmrFtSAhAvCpIFW6jSbBgu6RXmn5b3+m
mT0HYeGtYuwI+0U4B8qmnKU7HjHt0jqjkc779LIg+dyJWXM4Rr1DWW+VcIj5ApU4kIPnB5VfnQPn
B03+NpKTmtjoU0T7wLyyw4tFzB0iXSSJV3jeXbHtSsCtlcmLoBinHUv5zp2xbRiuymxGjWgFjqsa
gutgEBiosu5qlMOjhBBc7/YbmOPVjvVnruyTrc/EvwWPBIetJaXyY/7a0vQsrjCIuEWyGw1jobwb
xW0pz1svjhiqftncXbnveXXt2Ucv06o3HVbObJhLzKktcYmJV+YfKjkmREsMjxwl2+rhwjLsugKD
mKCczXe6khm9DZZTmgps0SEEsoJLThS+XmOfjNx/HbrZpEE4qwOCt2NgcL42AR/AhBuK8mi6Ly2/
tZsQw48EuPh3xkT6RT3846QkrLIgNOqpVTLZRXL/RioQ4TA6Ei0717f4EaGsyJUG/0zYDwLCx78F
lmSosI2FWUJjTiGoe1T04fZzzZnh90saKBBxoR4Z8DZDOubvl58xPc/tpFm1O4IXTQ+zYtrbQmy/
C/o9sTW2nTLhgVe60F1NoUmtIudofsgUXMkED4GeeKgG9g8vWuoP5BabIHLmiBpOAjqFKxu0jGwX
zmweoDviwliXvabSEVsMrKKqdIJRNa/irzvrEKlZAdqTx7GvXsauDbNJVUkTywISaDHNOgyXd4TI
kHpH48KVkyq+NgJjP6x9xzMsK6wDkV6xNlbiFvI/6mlq1n0Lrqur8qFwBX4Ja4vHD9Mq0ZZzMU5j
a1N+91g137by1BfRapWb2SYhgQGwKMd9m5lZrwmKzHo1leWc1diS+oTimx0rATBYR8txmR7qgJyp
IezVBFEimzCbBMDZajLop3QSEJDl0ThPXEG/N7hCE7B0MVsh3tU/SrwbLOx4e7MrffegkhmHGgt/
8VX+NCc9WLkcD+DT112o5Fkvxx0lxgNnf7xS3GpAz34RvkbrrKeg9Bz8KeNhRn9CezP6ObJ88ET0
BI8ILDq796jIj+iJ0PlE4aKjYRSprFCvvnjOHsZeUDFLbLrpwzCB8POebosJneQ/9JhhGw/ATqUw
/48aj8LbwZMBBqg5X1wVt0D4EXi9F6lRBbmzhLlBcETYJqjXtMHM+RuvvCHUSdqugrURF6J4/9jH
uOeWg9HTx4HUCqTcx1q1FgqRP8pbzZnAVobwfFq5flsV4AYJoebY/bQQ73Q1sgW08HRAepbkeVBK
okonk3NHMReCQgyb3l0dj54X43bZu5pKcwBVX/L1WYc9c4MLcJ6TJQaOPCOCSPQLNwSKvH19isKz
OotpIOO/b6AFOywbuLn24p0nP2OQLty9iyU7Uj3twYxjemevCIPE6Y7BWLpeTQfUzbGt5xsEsbFb
fHq3fnHU8rjNmkgO6zkBWcrCBhSoPy4Npqi4fWCIaREtRRvGiR8oKkVtxKvW7W00s+F9tPN0r2o7
0YK1z+cQFFJU08k0Gopx5ufPhGhC15B2hFemFEVOsHQXkC5qIherTNVb4tWtCqfsnPUCS44DnW0t
w0PrNgf6mUGpZVTdWVVnVDHmsq/mtfj5NyCpSCDpIaDOZ7uRA3TmksqfvpjZxVgaUUOoDpe6EcGs
vX/2v7o8SmPRQUmXmvl847QMPVK3gBnLEDVUaOIcOn1JTDfgdwhNdmytnggTz74iwNPgFucYgDUq
ov7gdUppyGjebEn8nriVqQclNUUJGpWXw/UU48qnAF3TlOyg5nt6dLPePCtfG+ikgrFnBmsPlxaC
HMPDHkCiBeAhrXfcYwIBG8nIFpuTXc/ESSP3FJJWIZZUM8qjK2ttzVVg8zySOhqXrQL5ajIf3x5V
RXdCJoSPoEF3vbqb6WGeq0j/t8Ii7PG5oulFbjmPTL3WmG3VxVsVvfY9CE8mW5I4pPNd26ZVLhZm
ukdws6yfHFvYaRjwXhifRdYeVMe1FXO82HEqCfnUsiRLViZMVd7glTbDA/z2StHXBdP3QMjIQZ0k
tJFJmqqzd6G1GNoJ8sjRG7HQhgqMp9ZmmdmVrl3Rfhl5WrrwdfVod50nIWs9obmz/j/9h71Xar0F
5Bqthb+6/eCu8MrI110pqI9G6cDjG7T9C4ltDSa04yEIJPFvAfdf288z8oy/wHm6cB84jXLO8KMy
hbSlTNQdfPH29M7/OkJ+p8FRcIhdUD2q9K1Q1I+6lqbit/cTVULZEeWYpDSbtw1reuZ1qO4O3UYJ
DBH5xBPtivfzHA57unI5nbY+PgTt9iuSqFUcEo+Ko7qYPvGk/xMVptsZNeeHqea02J8pj2PsDGw5
Zcx+P8mO4Wpw3zT7PcNU8ZbN98rpcjppsG/IH3G1z5/Xo49upwNs2VlT18hXMlPntvsNHycQbwA6
MAVuwdtnoB+bNNj11lq4HA6aQ3YIExt1X/MO1c3dbxdpoumxj6f/ZZ2ifvOzdiiBApWXd7gQZk/r
xJYCsWsWubLnzA7wrP3W8J4j4peLU+NPH90039l+pqIWnMWJYLgcmjYVsSweON2cCrOhjl2GFe+0
3Ww9hjRieO7Z2ipcMcKPoTgMgipr4u9w0B/PFgeOaARrD1jl6ah2r7OJ36jPzl8Oz4SQnvR4dSi0
gU2O3ero8KZoXr12aWU/+yXvh6Ac+IVtQRUe1AhZebIx86p9ojRNcWyROG3QRpaAQAX9jOTvj6lL
jbIE6GY0auaKkgNoTxxvoSMOHZEWW8+/tmmRRkcGVKkOvitkV3hk7uFCfN0LNrsLKrKoboSu0ioX
tXMsvRcbK8Vmd4T2AsWSJkzdklUI+wttGA8qEBaJSUTNynqlA+q5r9yKJjCh0vuJd8Vl/yCejJ+g
RYta8wx3Xev2dBUQkIFwAUCcTwFblsMEbZqjSynHD9m7jq3yJ6XcPov+11UOwIQHbObrT13YDKnX
RPc77mUnde0BriaCPm3KvBMqFFAATN5K/XP4uNhxY07NwiDBviomquasceZKxWCARks1/HOeo3d+
nIlzgkQGoRerWCPGHMsazX7AERaR0GkIIgeE2SYIigkpouU/npc1Jv9gchEX83Ckdr/yD+8all6h
cBoUSZRtWDb/eHXcKUyUNo5E4M2FkpiAk4woBaBVwatxURUR3+hU+aDPfRvQwgDtivowjEfK+Bp4
CbVHBMmtQHt7Ydg0J9XBEzFJptRFLu49xP65QJF/nL5m3mczJVxdn0VXuSdGvqEGexKlHlrhAuUx
ZDfDS7Y7VNc7zejDNTLOxK7ouWuXy7hvDWf0Oi8Eq4ZGDgbSLruytiw1qZQ+IwL1f9xrIWxTcXs5
PpeSgt5j2CYxWAq/mGSPk/i+AcsZSSeV0UL57aKptsCfaudjbay0o+Z0W/PF4ihfo1Q6384o+NKR
pQPg/1Y8MLPSYfw79dbV/VwOtsuf68Qjr38mhxXtbmzk+vGIV3RiGuSETV/Y3tx/sME+Ix3S0KWI
YH6g9ojsi5aIIAjVd72Tes+iXs6XychYyLx+BhILwPi4GDdYCDRQ8/o69lX0PsIt9XbETI6YUESL
FwITURarXWS+6bbBnbo5i1lMHro3CAMEcXZ5YD+on3pPakcl2Im/AlnJsCrXKEcoDb0/JV+io6a6
xgIlrZVGE0g/y1FeKGLJdmF/fPIj6abKvBNTCF/Bu04/RegYTI02edKPQdcx8eZaGzKSdQ2NhKKl
relCtr1M07/7ygcMknNw5/0k8M8DvhSSD8NXeHhnCZ1MCkqcjDjZUSpqjEn+cnoT8bpiejoSFdxS
A7NLkCyAgWM0idBigH8mCz8zjkIkrFNapb3udkJVt+oyHZrSR0q0+PupoSh8Iwtjo+f8Uo19bIaN
kwrEDekpLKN/rF5GLgbbwKuJWvDQa3o7A3dikJyPvJNaAgCl/kod96o3BuQN8oDUstl4PzbgvqPT
YfXlj0E1QYpy3M8Sn5gm9yQEU63efW7XHigOEsf2OGmgdbQvrtK7OGmZS1sGwrbVsQDeMdWIQUdr
/BKt/GjEeXo6lripZiOC8lUxRoYJC+R8IwI9g9sgetj55LvXwBRcgIh/TgQoKtJ5vvanD+k1FO6a
8g4i1NjTQ7tQdwED2eCA55hfx3LCxU4hvoVMqL0jd1nUCYDj0m/BSJ1s0FfIPxbKaNpdWQbW3dno
MD2wrhpUSX7oQtLPBJ9G91X52JSADv9nY4elkyijWebpkQJWXR7yh7SvqWUcO9gE1ytq5Km5Y6+G
lkDAE8Qy0nrhyMDzzBs1dieKGkDSU4GQwkePsJ8YaYCAsSvU5/FDS1Apkll9dtEy2YJjmDQXRy81
X6t5eTgiJaEqDeXqHBtvPTOBaIfjqJ7ID/x7sQC1AeSf7djCHjwHFH4zAgMgiNGPtsx6FlhcW+Qn
n2rJrRhoWlnQFigFPSmfs6HLjBfdOBlrbvsGX7Egxg8P38ilq8Nm6FV0cE1HUVPt6imKLrmztBI0
jV/zLQo3grhjursIdkbO/LlWVodkuOd4lU7BQCziRWcDID67/U5aIo45x+iwQ50p07eT+Egeeeoz
GiGAafHty84RbRdnEowW9PJzYeIJ3NP/SXCR4VfIL8Mw9YkR/d4cS+qkbLfbZnufoQxqjcsuDg6K
iySDCgXvrtXE4XzpGyTv89peelqL5pGZqXgYRLt5k+loLPKBkPSl4SDHib5oZ1dKf7AuJlTP3Ky8
hz6tfIgzQpPIbbzS8Jy0vm29CV/J119+2BKdj31AjzsM18xwYo2tzKs3KA/52VmVoPwLuhjbWLzE
eBx4Au7e4idQiw9ipnKBp3ETgHAg6wZQwld8BVdgH14s79E0XHQeyzeH+JkLeUBv8WMnTbpwbYHn
B8lvp0l0KJf451RMhJw+0f8bZc3zKEltsOJ6fUaeLRizrL6NGojdI3qQsltUePZmqRIO5B27T+jc
tpoN2l5f+7+xa8Y4IcXIMjhYgXDlJaTp9wD8CZFPftUl35go17M6ZtYpOda4A2/DCvbzWUHw9IBv
rmXN5ni5a83fBTlT0Y4/xnLhfwGfmvw1nX11Hp5X+/stbks11a/c0gUd9rADTFnskrgi0idaW4lw
M6a5HC3QNPMaPo3INRtDI7kix5r3QgNOTz2SIh9fG7o0O0oAYCK0M/+WxrkY/1aMkIe7bFupqKt5
+qC70BgfOBPV1qNn2XV8xWw8wXyE9cjyZj2lKEJ5hxvUqw0olYk4WCqMyi9Jl1vvWdI8x4wvvKlL
JKlLEZ+DkKZS3FcQ9rKuJABC9o2X3d+XbSBO2DGzgWVzhQnnHRYQxcKTACZ3GeaygtXOpnqsu31q
zH4BaSiCs6HkOeME/uiC763wLsLTOuO8UdmqbeaI39PU16GqiZjdNxEkvFaR0D+9yb3s3ggYy4LN
ozb+GtDfWpcvmfz0OGXsigGUkESehUqOoLdCNaNaj/fkm6zEhoDeQPOK2OP76vszDzgYDeSk/AHN
YPyAzi3b7QoeQxO+1YCacOLMnX2vBMDryfAY0uW5x90o8nnUw4BcNyatoGTFo26CE3jN/Kzw+e+f
V3bkz8MCotnUl0mBH/j9dlLjNC7HCoKKMJIwTXOuEvCFgVQN0aM8icuJZAjDIj8qEP4EuV6+QR+g
wP1uHNTTf9lAV8saiI5yF+shwteuclpuGkWodVTugiKQ/3SMcOXKrWPvHZ9MFBCejFwaLhXU34HM
dYa78s2+gQkCqtSLjP2tskC6RhcPkOuojrK2hMzuzcffgTdq5h+Pq2sqdlZAPUqDBTH+sNAXQKTQ
1X7kr1hXQUD0fhtRBixgvhaLl3IYSBDZxautI9J9YrOLaHMBNvmnruAcT/zK+0oPmGU7BoYhmyoq
addV6nw1IMYbjNboO/ItIhl6T54GMpUddGlP7/Szp7fJ1ZSFrA4XaWP/uGBuWg7NFWZf5v50j1Yd
eWW3o7rfKrp2RIF0GUPvoh4bZW0+SMeLKdOaB7Yr7xiU6N42f8v0k9Y90Oprj3q/s78mQRmMfD4c
+nCYWqaOwutfdd3U+ffuzV9Izk9+ilOZfHhtam9TFUU6g0IlbAFOz92thpMGMuM2zaH8FVGXgIqz
pe+ScvT8rPhWhUSyfLhKbopH4DW3dJPWYnc07FlgKwm8fl+m7ZfIMsZFd2Nhf2oDqXww0+ol1OGb
dz4rZfsT3yL2l8oT8IIW+mfVAANgadmwXg0K6wFdhbYVripmMDZ0cKUd+fLG682xV5wJKymD8qDs
3LexIyuj+HoExH176sC5aehxvTFVRcrIYQe0JdMPGE/AuxRVQDQl2afGaTNaR4lXRwE8GHIi3QQy
KTBF3MlFkgYHsDockg+mEWe+Yk9zHzurbpjdgvpgFjEP4GgdqOHitsXAP9IcwzMONMXTNU8r4IaJ
JPF99ggh1QmpBixNSlyc7ptANZDLyjlhHCX639HDhF1VqDQyXTRG4sbbzsznl2pkgNZB6+iVgyqq
RGCl1iu61wBwwb1H2vtpb++SaOZSYvJ+W9k+h4iW9LlJjH4fZ5s5yettEy495Pm7XLlzXizIi8cw
A5G26s/XExvhjtI5EnkvLNpXQVpbS5TMy4jHAnakh9pmJ1JWbR4k4j8PgFG7/vfrCGYK1RRspqhF
ywv0LNbNEpyagVWoTPk2UfwmzrXONvpCKhN19Mhix/OHG61xM8wrVGLG/qq9wfVgDG6qeAbrIZfA
SbCx4J57F5tXrWu6osdsSKhipILiNAe1bdjSFZo2QbvCZdYbVeMVOZCu/Pw83UFuuMsjsNDmH5Qt
VhiE/ptlxJXvFp9T90n98EGMRtoZe6wDYpikZdHAH90+rYf2FZbrdTEQCotPmpn3eytdmzvnyuoE
NKYJnet3vAgP6/4HOjZwzB3u0cycA3jauWCJF3cD/uJwirK1aVmHS8q09G9Lw2Hor94/JsCm2Smy
KYcWyDGWacTThtG1WU/sKIBsafUNfGXrKvUiY4rYbLUFG4DJVHGjvaiCDN5twhcCGmNSZww7X2iS
AVUrorA7sRLcxaiig4/EdIgGMHymJcv0xCulOzy+253F5mCPpW2UJS+Sy/ja2hZNMA1HNFTTX50S
KK66jN0lLhL7BZoLhZN2jENS1woi40Tf0SFCoYRK5+uBIEEXFUPES+V28HJWH0eBWNQb+PD/2ii5
B20BpvNwZyODXnB66kvzQBAU3Mcb+BkWkugf99OkB5A7UMPIC5/qFr4Z7I7mdXPUIMI4FWWnA2XG
G7iBIL/C/vHBXwP11vueaGBoV3jIMCwnr71HUP329H6OCHAXXH3ddyxb3dRytevZeK6gre5zOQMx
+JRubpteHYvzDJGdSHftD9a58eoH0LE6Kf1WZTJ/pVrMtQuz/AEaxFR6nstTJkixggLq2RPuX8Wm
ebsvz7rCi/O8moY5Wn/TUs7w2NjMRgbu63HpqqB7rQayLi+LXigQUSOKlgxaknJLh1KkyA0LHrdD
hoSn2ISMjuT6+i1KADzWYe0DYKkpudlMm00GBTaIRvG4jP16NUzaIt6lw9KoXgWpyed2xsnS5O4N
TfalzxAysbTIRZnUoMuVdFA+GoZGp0U7Zau2NetZr4vYpUAJ1EA91gydDLpCJu5Dhb+zWaEtAQJ9
pFuSLNmiAyE+BXoTzKm4eA1wtJElBjDpdHXS1GybEKAe3jL1XfCVaVcoPwVGEihalNwriDRXqjWJ
hHGEyojludB9Vl3CFPetN8t8B/7hNE6J4KbS+wzOKiAQrV+izFFHRz0XQEj9nA61vOA9+9x1l9Gc
lRfn6bxcPBhjSHCCktqqlrCkm+G+KDAQ/h2/xTTdqYi1svZLSJ6y5e7t7Cq8aW+INkX2B6VaB7xF
0bKXeFKwlqBr3gbLiv1clcnEiU3yKM5Bbv/ESnrMOq55yA6zlot6mejXpFhdSoutxyZgHm5K3SfX
IGP9eDEw4qW5KQGjzF8BnDxHDg6vadG7o2g1L4AvMu2eYtzata9PBrLDLrAYkqHLHNgpckAKgdUW
Z1hW4Ly2/Cuw7WC11ygXYPrKdvKiyXS6lgF+5L8GBUpbxStfZWin38k+7hlY8e0sRHY7f8spmYrK
LxuQpXnfHLwigWeppV3jpdxucylsbqWnieEfpVTNcsgwV3quHgLLfVzl67NVRGbadptsQ/lnI6mW
KoNaq1KpmhfBDXDw5V/z78int0dkv6njSdBstU7ZUIEmgnpT2JkglDoFI0rOUXyNyeNbQ6dp6WMu
cPi2sw97oBIfzdyz1Vus5zHo5I6ioI2VrmZV2KaM05ef99aKwtXPz1ZMVuKzHEZlZ9yUANtzFPZl
dT5RsMfQZ2y1ei5qKVYpioWTuryBSD5DNjbR+XiIXq4i3H951SOaahHzjMm1NobEWsB5uRXERZPk
yXujdOPI8Kyf12N91pkUNnKdP1bhs9AbTxDNLdJ5lQFaMIVP4wgPMeemrfmQWr9kngAIR9TvJHMw
KiGGDLy/7Mj+79rAep3qActObyNkP85ZiYSLoPSb7EMtNhTsnafvduccxGx+Tm1FUOgxMLA9jWfT
Nl54O/uSO3t4fiUdr4d3X9gtz2FZWjxDssq+FnHHp4nLpOYC3pTV25OFgC0yzInw6Wiyz/0nTeYK
mMLICr8lF5bf2LNj86Wrf3Q5pg4uJwpK1wLiKWAEKY7le31yQdJS4oV55z5GSS3nf4XMFSciDjE3
Vu5qGqPpHiDhELLaYNQCFAE1wCPgNqjAnvTxNhW10OwLGPCJmtFb3OhWP3rZXxulbMrsmTUYh4i+
L9x6XF7oEoc37vaFeTDL5msTNkgKO4EKRPTr9P3U06XZ4Al9TPjX5alG8rPGMJfm6tfF1Nd4rAfe
GnWTZOaqa0D8eIicdhFbeca/Ol3jwxNIqQvROm0i/4Q+YX1btNDAjxCJ1D6/RApH+g1+cid51wb9
71Bj+lEwMYWuYh6kMe8wTkHH4KBBWfAGbEfYW+VtIpRsaMqMl4yWRCS7Kp6nnGbsZDjD2yTKrEI7
mTvR0ucxPE2aJj2veRBPoGNV6hZelF7DRtdqGSsz866JbfcRvdTkYEvbj5d+hnMzBFOTY1gV8Zjk
6/rLNZf0zDwlGcM1WD3juouxhTB3i8K6DkrkdZx0SaVnwtD0OBXnAC9G8IIUBeB5XXpOu1R0AWT1
2Qb+ZnNSFDJTGegSkRumo97t202cMBtJbzt7DjmTDaT3HsNLXiTHgm5EjF5sO6XgWrW2UU3SOM66
Uix62aKsJVCLsRwl/wn0oB0BlXiHUP1279GSEkAUOCiS8mBrpCaYWwICLOMe0PMl+7SKCJQygzlp
/S/LHzrJ+xhedf4X9FDADjd4bARzAxFSVx2LwPbLAA7Xdo0f3Omek8QnTzFttUd3kvAx75Avu0Xt
BhwiRiCBszujueGFykATQRlRduGIEVzpq1GryAXgPamspU2e00GpRIyt8cNwTCyO1hMLWBLVGW5J
wrjCcCyBYkKrIukBz+IRIVcCd9Sjs/DsS/yoPVMuVKxCL3cPafevJn5/p9FgdbxhMtCigfJ91c58
KKJanBI8QrGK/sXDQZp+ZGB9Gc/P3NMvuVqSkyjg0vXzdoYn0WTUrZYtw9Ubj5kCjjzmuiMiwuaF
paljcWEiWyluHnPdod1Uim2iX5+A2gX6sg8I6IZa+LGdoPvn5yqOg8PfQAwtIM/UaDiYu9v3uBi+
wy5+aaX3yQgr9s/gFkuW8Iv0agVhDubtTijWHjabxS6B2/MX4gG4CepFXsnoR+LKqFp6AuMQxn/L
hLTC1sIVqrtpr2pqQngyOHlEMO5oo9QNhLk95m8piBC8G1U+MxJ7DBs37BFrwzBeLQa821xxOEOV
69aLi8uKHfgjF24qN2hTK+rQfkXitpWktJkilrGEa3u6v1Ed1LhUol6qfImqUbLCHPnmtWLXqJ8w
8Qmk/SSQEFoAXQ0RVmv5PtUhaOTJcm2RzWoYaqivLZlvk1Mb4BvHASZKe5oiMS2FfGf7Z7TOAloK
BAgrSjV3IjnZEvdROMxBoJJHgS+Y+QRo356g9ZZnzqQTnmBWGXFDDY5xwkXqJNNSWq7gYmQ3Rcac
Q0O7Fu1DcVO3SEEiCBBZ2pi72m0TyOMgvoFiterfuiWgudLzktk49DnV2XZCbDOrAjhM242Rd6W3
kto1hiF5mCPjW1H26AzK1kwJSkraqQQ9kxaQDZu2T16rVYev8gBnXBDwNoY5QsnErjwxLuUJaE3Z
XMaeVqho0wm/pua3f+RMUM5jjD64PCoVQ8Z1XaUEFLJfd30acjUdTYidGuODpl523Oga13RIli2L
pzrrXFVQSQCn/Bt4IKzbadVzYD8C+rh9u3wnpimi2MdeERDHRtZ47ZJCbEMgqkRxmrS2jO5GGDvc
Gly3OnxvIEUIcESH/XbD/S2TP2xSp896kUEGSuO4fUKHvWikPNI3ujlJgFgX7dDL4c9f7KfOKzLa
OA9nRKmCJT97aRrAJi1zBJrRZaR9ElSXdWTyR85sDlkizCY8rQeWuqJ1DpdRCXFJw58jJbbdWMSh
bzCMkCcfuLPzHLv2QOIJubnyt11hKDm1JV8jHJSoeQrza2e+qTVLANmMNWuZKmC0civBdFjq+Nol
oa/Xn8+SF7IsflSKmiAoQo8sKdujzWBveJ7iT4IkOh1IfAsG9Y/tOX1c7pZUHcE1f3nCHj75gmdJ
FPPeg5p5MFlXUvMaromDAWis+xQZERrlYvasETUNjArNTkXKSF3j+8TlAh/8eJuu4UzVIZCcF3xK
jtJY10CGfTwo7oRqe3rgON9T5P+OpQFbbo1HHPPm1dqfHqqvCZTn1tL/7RG+8r/WZlzMRk8U6+nf
deIbLjGa/NyyUaqPndrU6z37Xaax7wpcsh5nJshJhuDjHQZiPmh8wfMNrUd+Mna1ys8dkGsjnXXS
tYXnD3fUaWCnp/koau4krgZwbASBBmJgi1zFtagPMpJdjYGLo4h+QzduCfCQPV8Z09NiDkeQWC0o
cyncT0mifWrkMyAp8wO+Lx/y9t4cOg1/UGnpYhUh1W1FzuAbFz+KE+R7+X5Lco5Y0vvo0Qga9kFf
oRwUsBewy2ZJ9OIgDnlUBn7tR2/+ZZaykqdXbJ7Xmw3puQPMEtBdiSGPrcqwgVGEYQC0dkcOfq2d
4IBeqzzWB3FnYomy6T+QnhKV/07aA/agLoQuMugFlnYkxnAcRRpHrF3QlgbIniwQqLHphMKE+e48
3FYMjD65iJIUOsQBtcvnytUgGXfZ5W7N4YUCKvlBwmIxJHPMfKSJkZSpibob+dDyI8dO3YdSa+Jo
m+OEgYEqOt0uImyTmsq8wjoP4hpoRiY8W1bpPJGtxr2RAgUxZBTG/w85SOUxrxQFWxmPPu4wkfxk
1kEuZ9adxsknhlg4dh4ki8vjAwdvYDG/ePqlkUvV2u2L6o8CbAC2mlwH0JAJmll0a2I728yFcr+E
7LLkpAN3dSXBZWjgTsB1CrU4vqzxJCVUfGu9Quiylda9GgXNLHMHn4eypnLyxrdhJG3v7LC2k2m0
Wk8YbOXGKW4JpH81LzVF35uM06tM9ntdFb1XZWGo8mDIY/sv4bVswk1c5+oDjKMSl0ZMTxSNvvrE
ByLABohfrMhVIaDsRTnJEvEyqSwABy1ZfYLlU0iyZRsjkVjK/53nyI5Ht/IRTQ24IDzdenzTV/SX
ZwryeFkMFi7J8MYzPoEEfAm0rHWfkEYQjsz1LXv2x9BSPMheHYaHOfI5Oa411cS6mWRBARtRZwFq
V+8oEuU/fOKaqL02TWE4eV5ZPMv94zKAOe94GhaFD6BlFCUHx9FQXWLqerDCRXdRdTzNyNb7kNaT
JQcEKLX0R1WkSZMYuptbe9GB7De26TIXVAWS/NDpu5qck2VLYjJrZ+F55Cx3fw0lCmBzU/enQkD8
x4aSTYySxWKOopaZTG6NgV1NslbQs8LHe1zF1TCDxAx6bnLOESVg3pkpA4yHXVwUyVKqNusiwijx
t4doBMh+lgK5XthI/mjLoKADHThM0yvJj/68Ss1CKIXy4UG3H8XlNUSHNbAwxEb4i6TUtN7O/wR0
fTe/Pm/z0/olIkaVy0keXOrNUS3mrJmMkNKx/DXiVDlAsnF2DjG/fKhzN1fLj+CxNfmTFX59mG6J
uh5SwCaDKWwlYHFv4VElK2wcjzxY+FO9sAnG+4SymZQPa9IPdVj8ti6DCpFggYsNio4Cw5+aIIFf
IOMR3dOoJUBVtynz4FQogOgLuNJ1jmj9GG9LyO5xgrHvJDYlzthmuYLjO0ojbxMx747lTEVuE9CW
18A+b+//Dt7wC8Yz/Byb1KSS0tUb9f77ThCdlHH7D4qHBHIYZMtbqveztslgC+0cOaQpF9ndBhJ1
rE/5SEqOGByxW7VY59gIHjj5dDkgyYA5Dp7N7tqw9ljIqQklqloSHeQ271xjFP7HorULT0ucw3bT
H52hufUoKeX4citwuIlwlT7LIPgnEDV/VA1FOufyG0+j87YZfLaX5rOomph8RwRyDp+fjaKYo07T
l9e7GOYNvigcyY9Kh52xyMc3kuHN2qg0KWps5d51fHg1Ry02v+gkFN7xnvriuCAZeR7OeBhrRmhq
O8o0jCG1DSfbMx10F+endeUtFjiq6eBjrfBX5/Ycatx/xZ5ijLe9Zm1Ke5A+yUOVGtu4LDS7V1sn
546l9cHfur4kGc6H5wmL1C/BoSPnOD9fOpkXsvz8GO4iDXsZBRN4XyluK/OnWWciygjf2qlKrKGt
ZL/SZywjpO2V46tXh4IU05s5bIIaR2VyG8Lkbub7YsKdtSEWpJ9XIGYyt8/H2LpJbAqUE2Le/e8t
5CSPSirPqo6CpNKxtnlsiy//uh81Rj+v8m8eZxKSXbgYpYQWA6VyWJLqNKOhA/zPSGkzv1S5N4jP
MP5DSBoQY5lndUCkICCB7liASZigj5vfvE14mAtjHATwMgs755XrvkAyy+k8crwa0vPR/0TUyP0o
ZawpmYHSyyCHRnBMpxIzQMKeF1TaqEXy5ErzAfFKm0KhsEE+ynBnqFARCKdIqQ3gbV0lnbRnPCi9
ewLbdqzG8oKLPza57zCsJs8+L33Dof1Q9gV6PKPyDMIBr6NuOcd0FdfKPzGjwowaBUo1Ls3gw+f2
5VNRbf/TXNwrHdS6miBnbMn47h2MYb2XdRoyU3DViWZrRb4AH4ceA5HpYF635kFb+lq2BKIyBuoI
PzPn58R/O07FbGfxer9Bb/7uBFwrUNRCSPczwKLOvoKPrvHK4Vvp3EfUTtC6Lmo3gV9NnJCiwZ16
8AAD2ETf4yA82ITC5isI3jUWGDPu/nc5VlETqcRtYihWf4i0X6pZuQD+EFtTFwE9OV2JGFTlyyk9
gapf18s1M6MpcqMuyRk+4MS8D3WuoOoS7yfdsuR5qhlPyeRWDlVo+qxWE9ywDXqRFADmS6oQ3v2S
ZW+euh/uQhcUE6qTj+/KuTRZ7J47Z9UllKNsCvnvcXwflQ3c6yUAroH5w5ZLROXHn6G++MwkiCbd
o3x8b8itM0EyhdPt+su+Q5/vI0ornpQo1GsZOQaUA0s/ShyGm7lRxFES9Wb+tyEVNw1cHx/0Gqxk
o5oX1PqZ2QUYrABWj4pT6CHL8941/d4dnx3nbMAr0BS0UvYKSZhPacEBfHOHERmNWE851otXASGL
x9sN49B8PMcR2HC+GDeaUVNHEhg2f9/XuI6B+IwFT09KnWtebAJ9ORGy4DsihzCrCPzopTsY2Ay3
TVFw5iRKK+BuXKqcOD2onETMGfk+eu9uXaBjkNvlkpVglbrunsz9jsy+qxV1BEBESmXLoemlou5k
OWtiWc26r4EMJFCCbTTSlKWEKYadmS+a0Ya3exKVuCTnu581sGpky/XPs2yYTqhsNrhGQhXT68oI
6DOnV7ynUjaKIRepkjnoPJ1JovK2tYYH92dhHOa++lW13hcuT1d9DaIMn48LrlhsNzS6A1CfZg9Q
Pr5+oLFS9FxcvBfctUBOgNBToiszapfnJwuZVr6ksf6llWHklZrtxEocaMBFXvzafK4KpoXU+aOC
3aUK2l9PWqN7AiAw+dN09A8qGxWa/8yyGbhQ3R82TY7Yes1keF+wxLLF6BKi1z2Alr2EU4In8FPd
CvuwTesm1eBnFMQnckTTAngMhsFR6FPGmVLkwd7wOilWbg7ium2W/AUaiyWJvGIXJ8pEVlW2beTc
T1KT6lm3msSLdpPYw1F2gfWAhS5NVKLBsp7paQU1ZbxhOrSvYd7QaXvK88rwusn2VhHEU38Or9D4
l2szt7zANLEyoTGWMlKDWPXDiiJPqEbwKr/0PovAfG3Bu8biea5RB0Zp+7tofQ0dJ57Z3gJsjpbF
z/GTdozakpI2mb7z2LohqXHQT7hvaGl4ApZlIxenTAo0X5zBTNJg4Li51i8ealF7F480h1E8aSPJ
qLCzOtjfyrXHvhrSOkUodTekEoCRmYwniaVKpXbIBDb3prvKt2z34jVFoNmnuJGhtdkTJ/nvLhTB
gQUKps0wk4rufrPPiXyP14LPXuYDhiKDVxJBB2f68EW/fef9+qVt+AAnnUwjabAXtJhH1u78jor8
j2SQ4Dk7GmD/RTbmry8mJzKr5MPxZqIwTfeTjCjcWLtKBklPkzBSAwk9+beQtolE3P5QEkkhtYNY
K91Qiy06j9SS4CkhvDvu/SKBz8ToYkopazj9nzd7tadGQTWg+r+SrUAw+YqZUjvSvTcQQDEahDw/
27L6H3NSbqUueHjNqMEFADaX05c08rfo9NqSB8jjCkTw0+si15h6TVAGbDuA/6FHcGThTtCbWclp
v0ULK2fzFIcKKX4tNr2mIjmR9z+8+qFZUeaRWGi8phsxetbOiSB8ysKY/KoFXKH5QhbK7OaSoR25
s4hKsm3lUQ9C2EQl1TslbNvQ97GBrqE9e06nKQD9EGdBF5lZ+eUaLFNYigXiMCrwYo6BdvqzVV0N
DOQwYhEd7e6pOA9c+iawvXPSSKKuiUjoRz+AWtKNZDYlJ4pXMEPwzUL/IHoOKXBvg5AoQggv7TFl
CEs6YPhXelHPZlTXhNiaNLVq98XT7HtSDZkPpROu1GhzlT9IE6WToMGasyZPJF7/rm/VRRoNmWoj
AAkDNXecLccwRnMaxTkl/E/poisIgeKKhjjH+bb5cmJ2w4ZnO7tTEPVMyqYBo/SstUNkYKKA4lAG
bAjlx28dORJ5OR7hu+7LByDdOm2+GG5t/bMK9O0G25J8/7K2rRvC2n3FHbZjsWzroUIDsD4+01qW
QHI3cX51tHY37Xse3LBFRVNtYecznv/SxWYDWPFTV8gqNc3NNuiJ7cH4DIxzovYqrxcn9A8fkYeo
OrleB88NmjuTQR4RWUt/f+LxkfpNQ/MI+Wwx7anEH36PiZ5ET6QPeiAD4QCmI1VKCUZpwVohvvsx
vq7fCspRQF7E6G1deI1oecc6onvh9zMKle2Nhz4kbHzRb+HJoMkhkGhyYoXiHZ4hShNRH6HTO+1r
c2Nyr/W6xWlF6eSTJGTuL7yr2gMJcCYxi1pL21RHy+ElXV4r6yZtDkQzkxbtdwvd/TgBIorvkL98
akAUcroCMu92+yQBjDq+iiSdMdY/7AHS3f/MZvO/O77z4ymTfiwGLZXn9dIRvrSQ7G7GWx29Zlyc
vskOPTkyXjqYd7ygJtvlbcQDSnRXXZDs8ZFpjcm5/uIpmYJmQ6XzK9rD0wHNa2UYhOCnw5c7lNX5
3Vwno1/edUfmhoTDpnfeg7GtZvDLmckRKLnUWCiN2LhD1oOeCnMZvQsz1kOFihMjqHmCv9HXZraY
ihemTInq4fMbYelPbOod0ZrsbQipFds7Ja3sWZJj/s5ln92QI4WKFvy8nkDADqmfJ4MWr37wz23V
cUczW+8q41JnO7HJfFmBqydBBVOI0+XGxL2gqq5WIhZbKBaOHqMBP7vi7kLFVvz1uXoUuBPjWsTp
0EurjuyrszaH2CAft9DSeUWovNTpg91Mx8hzq8ueTBwDFJzPyBRrjo5MXYCxxyJ9yF6wcvtLY0zI
+4s0SgQeEZyETfQPqJ1nEdpjO5VtJHBAPozWuydJ1G46uPPaOAIvau13BZWdDi/AOQ5u8trDNkQr
B5psZy/PkCmFzce6OZsAMmhsesias/qvyQGzdgL1bJM5MrchuzbvL3DX6sk+sYWpUedwdoT8bVX8
Mgg2i5S61m0tQBvivyS3hURsH1/Ztexf/V19ED6OVMfQvNbcOOqkxFDxdNmwjwKkbqzQYjt1ZXoQ
qIWtjak4cclcACjPIlsx3T7Wy2sYZU6TKwZJgdD3eKAKu7p2mKeY/t2CdZ3etxiVWrx04kwCpnMb
8dJw6lHPBn7/Qbw2dt2evoqfPGEdAg9Pkyc/T462SbrQ+7gmHImMwRcBG1MoB47jUp3HINmIMrOq
VjMalSu9za93IRtKogdPM68ZzI3qjWQ25qEt2HTmUUT6wT3k4WtVRoF5pL6vrWSdnljGF4YwIZTv
wJBXEzghziIpKvdl/IJY5HZwF3qE6yl4ELIJVhkzkJ9S8p/ZHw2PfIJ/DSfBJqL50ls9wA5iZam1
+WltJEwghUoX9GoxjtrRfALM+o6paeVEbqDFMD96NF7JicwC/1Rebm2pL5REfCcDbPAOKNPkIJe6
3U+HS6/TvI/Cp95P7zD1+bkA8euEPdMKjddeLxyF8ETQDW8H8hP/i2QeTKxBn35bQAlNADrAnQ6R
ATMwt2l8isExjgh3vZSBRSFUoxG0jOud7wt4s42uv1LhuxxT+02eFrc4VeQfYNj0ZV5VnNbJiMe9
mxxKIlrNESJh1y15HIwQlWr1yMpIfkjn/RR5T2/CWBwlFeDz3oMKIl+FSBbMvBJG2rKLx8aRNWuE
mT/DbCEggqPI1Kcb2qBzy6pq90EnEA7MSQDC2ZTV6P5cWccyNupsTV0+iAhepIx0SFbEVoK7zxrk
RWthJKF4urz58UYWCcZgPyY6sqlhjh4upsDlnMtiiI8vp1c8j2lQzs2tcMlHv4k/zH74sbXOh94d
CTAWW05FnZQRxmHLUIn31WVsz51o9VLRc7nEVdYizoXk0VHwqsPV8lv5y9+fVJcD4198K82PyPNG
2ztbMNMsRxZLkOAazDAQeeQDeoUDYHGJaZyuKnMtmJ+rRIx4olxGduLNNhYmfizRAhE7RrXb8qs8
IBSYSgZUpmsz/LETXoWblGV/Vdj3DCWSpYMtP/Bn9GQ8S3P2y9wOZZAEM7aMA3bdmNNoQOm4mMS9
9wyIAvqVlF4sJPAWyGUUDDWJW0bn9VNCRQeB3K3/8fmJs4OuCe885ndb5ACMrI4Xs2TaJR/53h0P
PvlqKr3iTj+sGvYmd0sT0G+nCt6SuuOhM89kknUvLHn7MbH7BpHeR9xVNWEbYi0gz7Bh02I6ZTAm
DYqB9pn5cfhTlMKC7ga4Vm+nJSLOCdcns65yruh+6oIb5hpZ4SSjOJjvd4eLDLllJr6I+KWhZ8mZ
t6Zz2crdn8981nIHeHFXQH+l6oWo8h3Y12jip2/2zvNhkrsIQ2rpXAxCfbdR/kOTTTstCnG7EClb
0tbsd8U/qRtmg6f/s7j/z7Mpg1onl/ERnhE0KrBDRIP37EHXwpu12ZVItwKGp5xyDazVN82DluO7
IWoqJvrkzUgujwPiaJNAqI1kmqBR6Di+vR4MXnD7EXMu9gV6oOu9XfZgVtsWMz+byQGeS4OACWgy
OhOlYGw9qDKdzfV7zKz7RGoJJFFGo13U3dQSvygy+5+VFrVay2z64lWPURShqwnpK3kTO9EF1WI2
JFGoP1iAmuCzQ5pyroNXqtiZ1X56GY07m2fp/Nd4uQd1/6Ya8PXcL6bnZNDjvMVzzVcs/HD3mTbr
TWYfEpba3cDp4IZXnjEgufrsMH/mK0KZT51VIltGH9dyVskBgqKYFrQWgWJfkRImLsm8tBj8aZE5
YiN7p4NBdPemL+3v+eZlbrbMzA9g6AZmFBJfIax7qs9WiLI/j3Hj3N80UKf1pGW24rdwrq5sDPY3
HCQyhWq9slcIQEChxiXgzqRjolYhI1LGKMlAaemChe4TMsFU7ErDmpj+Mp3aERtVdRhA1GDptKBV
2rUyIrvH75mh2CVwyTvtGIBa7Wr2ywvOfEiFE0msIhkDxGiCwbfxJrSoE2sWBy4Fz8j3sQ31NXI0
O6ED+Tf9qNdo1JXZTa9kIebnaHSN1jYaDB1h7hrdr4MbA63XSEBGjOAMZhP756MbxAoGARi9W78a
ZDt8OupbCEOsWpRArxDNECAyEMuOdyduf7gTix5FfGRZbXv9xMYElLef7pVC/Yu4Sk69S2Mnk6Z1
ujnuL98ZwgQ4etK8Io/70hfl/KN5HDSf/wmjyDcUZGTHW+kcxf/m9QFcBpbuab3FoO+iAueg3KGk
24ZEwvEvaGgnWg8k9SaVznZBuddQFD8gflAn8vAUumgHw14OYPxQ92tqfDeaoNDyM08UJNB+xHKg
vVc04eoA0Wyc3j08PXHVe2aAgwNYQ5zo3nZQfcZhLOxqzmMdQYFN3Qd9fBlA4ExvIOVvqKP8NH4W
f9D5AGjtIp598MKHAsOdovJkIFpYCtgZCCRNvPRfvja+bIUbF39eX+2Ts6aI8ucoF5osJPqx2GZ8
o54juK03J2XI31usBF5j5tBS83Rtg5t4jn/0ckPldWN0wqUqHq2kxxWCJJT1giNmPGoik+dAr1ei
CxbA8oEOc9cOTLDz3DqrPFFuKgxH4FChU8OFdWnGE9Tc9BDWg7tpR3IXP2fv7W/h2/+QNzSOgLA1
9p9Fhp1EhZ/b6eLT169Kat2+cxj8WxoBMoMi1lwy+OsVQTwcMQAM+5sn3/ETNjO48UfHf5YHVDRx
Ap/axmDu+Vj53jwZV1stGasSDHHsCQ3au8199A0n1FuzJD2Yr/pG5XOEiNtE1wUgPtbZuAKwV7AL
baIdgfSCqvQQLFbBp4GlE3axFIwVMwNYfRaggzPqJyr2Bi6DegxFE2+oQO788aSk2/Gb/gtfwmBn
NXorJioK87EewbBxoYfsWXZV4g1sYssTJSI1LCt+TKkIH3pNGwlAME2rum0MSM9Kdev/FblXlEbQ
Q46303C5/L55GuTsaWdtpy5KMwOtbltMAe50QCETmndP4BGWmnxQQRTsCVnJiY7dXziBOXoigM6x
qPCl5OXOGYYXQ6Uk4zxxVG3LSpLEaAMlbqTOckDzj2acHuT6ddLxXdDSox5nk5lpoENhmQDXt5nL
qP/cnpBcmA0SO6vERzYtdIL0MEecfySpa/ZhnIpOiKhK3fX+TcnncqZwAeioumhbu6IsUZKMEAz3
hb/ven6z8ga7AdzwUCIOKdq0/0t15GO5+cJceUmupn2mLD92wW1pcfmhC4dVHhsBcwG0jv8OKioV
I6k0w2julFQi1Xk8CqAdMEzvo1jHtfFq1Ni4YVG4HwVk5D6nd3QdKYJXqMKg8BkWZjno0ZG7OIOg
bG0T4UnZ/kfF23RsptHoy9ZvNwB/hU3insM94Yjy3NLgm0jSPO3BaxlDWe9lGI2dOwblFZnGVKp4
GZLuLcSH8BQAEPqMyHxbsWBjXwqnGiT35X7NOXl8c4Z1BuAneguTH7F/xdNW6iX93EHFM5Rvp8NM
hh/EWIUS4UZkpcTkaHoJgecjqaiJ6dyHReXXqdgTk8inq+tkLw9QGvmuqxTH+pzr7rhZN2WmFpu7
G135mpy8ffliAbefGubIavFFDgcQ7RUYCxM7INUiHTacmOmeVt7ieTJkDnuKV13wxsHTi9t3qeqc
Uheumi1/cEv8xQcNcsAssKrK1ipECmK8ymRNu/9G0ynhIOu59oq79iXfERLH2cLo9FK50Ywp4Yod
EdV7crmYVlw+RE8XDzz+GRv5AH+Vt008QKd+MiR8xxG/NNrO2V+ZAF1zb0ZET97b+wXFwqxcu9gG
c6Y5aFuY/8PIIdiqqxvpzSH3kvNJeNY0wETzOAhHWJctox8k9m4hpwyjzxN8XmMxMjX6d3Al7YG0
GPSV1czbzCyEIWSgqCSPwOVuTGnkWWFpavxH7+ougK3oLQf6FGNgOVRw5pz1ddzXQ6YhQji3GE8C
mC48FZ4Bj8UD5SI54M94gjr8437r7cqSM1q32gQgYCoorwWMeawuT4SiY/cvTD9o26tHWxWbJUor
HXT9I6mntnr0WbxQo4rBW2WUHFNaTb2bAkF3ORxf0o1rloJtU+zboabJ9yG1VAnEJ1XqKd02cqaN
aANOcJ+XWam6fcER+UFK1ZmzFdOIz/avIuj1faAwcalQkzxnym7b5lzY3xeYVuiAZFofOcfRXajw
bjEELvo7cvZ/pUZLpsBcz1bI0GmINRBg1Dg5UnNH41g5y7Kryt037nc/j3ev7xMAbof5PWaYOB68
scrGrtAtTSMcSzEcpVFD9exzzJrrBWHwCHJO88HUAwM/dpsmY028TFJ9yYPG3C7Rz7/QkFVGEOk6
U5pmaCF1dNEBULsZvtZzi6IRQJTmguEFPMbfMhN+R7Lk1zwueUWycxqBSDFPFg4AipgCXM+Zn05H
1M7GAk76md172fE/u5ZgMOFf/XJaC7OlCfPB/MMKp+cfiCWqkHTdLSaJqdYFkHUi3uLfv8FqC2s/
lVBP/V3z/UVn5vYmM5Fbo6vJBogqXgSFVOC/AnDwszR4Ml0KNtUlwOuVgSOKOM8XubPayAJhdhFx
Sn/mfrG7Ew4gpyx/Col1bwc62Ed4OjyfzK7k61DOs4LOPOacmGkqJ8psR6PR0CLGwy7Jqnx7RYgr
qwp6cK84gAU3jBHlCW/AvSpTNla2L+p0+P6eMRIkTmCVuqkQt6YXXMujO7bMd+THYIE9vI812hW+
XUDjMAIxIIzazDn/lnuxxfDIDY8STfx9bSU8avahHOHfw/Af6NFmin0h/YUtcJrKMNcAK/2Ch29g
+eY9B33JGjVzpR8SaMp44yyUA2IguQVIm+ITQN/y7prZlXuFJiSFRqRlGFlqE1f76kMsbIJp1O0r
AE4ySBO4LAqDH3nVzEPCCpMFqdxHQoP3Oo9NEUhufTsvuGpKi1gQlZj6dPDPS0CH6Br9vcPLTvJ1
pXZFPXTBYBWfD/3wbmmqd/evOdpuge00OvexPUELPdniyHvmXtJStweHqMLd4oAyHN5587KuNWih
bR/fAKypCXnmPoLWLG8V1An+TknmSYN1RYileV6dT/VAbLHlz7p2DZMAx6mLtuwFQUMugObiCBWB
qMiBnz/uBS0JdqPGEU1bhgdF1KdDmmAzxq/sO37wE0fEMGyNvVD2nxM+2Pubtdy6ewqCieOTPDi+
R/kXwKaOzrFH2lplJSa2Xy1Nn6VLsPvcgEM+1gFC/J4xUyPZWQiktcUs6NUjO59mNTXKZTrge31G
Fa6dLXr+68tXyUC4o4ViiPh1CAhOBTO5lc7G60s59BzIZjcX9Zec3ATAmBgm1VAmp6+RKK0AVdFm
uA9trLvC5M5dcTdwOZxWn9fbhAgVXadhAqDGNQFiho6V3fRJHY5BMD0+vvDopVC+q1mPnpCKpvLX
1/grcpTLQRFooG8dNHXzPvM+RPuRYOnvKTFVdTHXiDN351LuXKRE9D5osjhuTL+ermPt97DTnhIO
xuHh2LVha9USqaVvTrwHrg7cc7sNxpvANeGTqja7AxdZijNYdQbIsuGMSFZcqHRm/h4wnJHvppe/
YFU/QhiPV1Lpk0Vnhd7EOv8BdoWAVaYaGJoOmXHtDET/0j+ML7D0tV2Z8s8Oj8Hwe9woaoUN4dwh
AQU/Qs0a4o0X+KpxUnuEciiQONwfvGHNv7AorS6ppnCZrCGFqcFWbJYOgDkGUD/CzTsNW0q0iBw8
tIIOqwfLn8at29v8PsOxvTqTssiVXLd9rI4XoK4qjmLT9OaetgWkBFNMqB6OTGAju5uqocAuoEXe
Tvurq1VKEDvoiB7H50zKJQpFbCEvyBlz0bQPlETc8KIp7vSlivbKchNIFTx52pBDtrR9BUFEx2de
xDlSYKwhhR2HcMhsTmqJJkvfeLoRy5N2B9VLMuGQj+8cjpUMFU1An3Wd+h3wOiAYBPDRyCdDa83Y
+laFf+Ri9X3g/QNW7pAIJoo6/kqK1qe1VXvLITkAJAkJUQAnwZYvbRoDfSpUdeO/fyzSnqogHknZ
sRtF5JzG/kwbhqMT0CP7ZCTB7oGu/chtVbFV+jlWH4OOC/vJL9apqZ2kVmAPv1lbqTPzcRutnQJZ
xOn+V1sW0bZ+EenG6/vHsix3jkpz69L88l2wCda9JOnVwjdPyClBFiX/uxqgqRzqIJ+4un2bd1Ye
0Ywj+TsGw2YHr+hxOLdjkl16hoJ0brc3dxMxfVTvLIR+lX+1Pwj3EtSmMDT59Oyey9LEOvzGiptB
PkPmte+dSs0JF+8YYC4inO85l0FhjMQKlzV+1mQ6np/sDo6AkUIb8fQ6iVeOqNe4yHMSjbmhWuor
EKfJQwRwnM9jzj8eg0Zx7JwnOtHSXo4vol/t8eRWp2Fc6BwYpsd87RsWcqrJa2YvMSLMWFUOwdBw
hpGU/bpB3H6xoLWB6IqCdRQZmwjDd7bL6wE7U602JB42fh5mLiQMKN6GsOaOe7uy5CwA9q/Ja1d4
DbB6c8nPGSeWfGs7vNh0zFamlKimgUc4VhKITQHkOmRgyRyG4jCaKpTcFjimMY1BCHXmz708SVhs
w982Ql1FMa75X4dNUxcSmWSiKWcWkexMtr00I9lU63kmuc+R4g//mIBgUVE7M6QrKHxDTRZiaTl6
DW88fMooxTtvegmCLjTUcjsJRTUyvc21Q6Sfy5MiOhB81+DxpChDQNJ9OCMB+f0hizRPg9a4ThCe
PCKQ6YqG8ec88SOONdw6+wJI5fuvPFDkkOVoXjbNYDtpCyHHCCuiDXfvHkwtRlWTSwOBkIspnK/G
gWbWRqLX7gtzwHZvea3oedRO0Xk6f+ms0NlcTc6stFXV9sc0NLjkQvSMi6mFozvRYe3ymV8ohJSf
/xuR4d0HRBF20vXgNGAF2mtf0c44LNUz/hs8Mlnd94oggoZlzSPN5WgcX3TtR3zNDhRTwEDcYQzo
SSRuCUrNNYLtCM1Qexi+G6RA37CY52JZY2+GB4ru4cbB1tuCV50B4U8daQkNfN6Tdem5B8lkscLT
wJrGDLvpVTEaGcidRJM4d4TCCRBlfcKAgQQz37Ye6kUXb4v6Cxartrn7IsWiGn5lK+UNoTZ/b58H
NA+oKE909pwrtIhSFdjnU27pv89GfKoGxj3vMTSX1YWnCaTYmh0015UH1rszdAhzWJ9REzhYWA8r
4rc7crEmdDMiGA/ST1A/bOUNkXqtFZWJGa8U8PWuLfWa0bhAvgFtk4ep1GMq3VLHALua04ggkepF
qdeiGsKQXuiH29m9bZhZWpPiujVg4vqOZo6bEDcLYNA5ty0M15XfG7yiG8I1F2DADLBG9XjjXGNr
4BUH67a5y6KDwPE7T/7z8lRaDPPGARrQYwfSm2+D3taR/LvHjpUkNUBGiDWaITsdobeLFJ51ssDG
5n/ANIaK8v67FEt6Supe2In6hA0rQRk3NSfdPT9FxOmKGOQUMDFMGxW2DeYsicAEj7r6iwR4Hdto
afK/05jaEeKlSmbWxLLL11h4iAyuYQtXErkqSDw4O4HHg+aDfCoHKGSbpN1dCQB0zxfbmhs99Xib
SfqYEF/HG4bB67ReHxerRJkSTn2MVLuhtlzXOGgJCFpuxGDvI+7shQBbtWvKrDs8oobUmmekUzQt
FL2EcLPaKA7LD2ZfNmkz9fPPLt4N5WGUZQYU7IjLLLmCFyUa/JgyLnMse1oiSEQzSsdd7TOP5VGG
Mlu4lns3DmUIaACAUxKwJXRIZqBNGE4zylahevFFppTsrHOuxwSE9axb9rmRf0/5VmmXs0xumGpr
P1fHRVSIUdCI4Vjind6IDqQEAcJNanAXBusV6A7T6avJVwxKVQeNQQNBs6ELpT52FamrQU8biZx6
+rVos3zgXwxURs9vuyxKwcEY/XufxN+sypKlrm2nxrg/kkLuf4KA8fmSpHBQFbBzWd6PCLbY22KA
C6fOakwJKu/FWkkjHoFiOLp4ENIyUg1D3ZwL3ewh+1MLjAyWcl6gNPkmTlQj5qKJrYLojHzFYcV/
65bdooxje664f/R5wpf5VvgsBtn5r4fdbv+C8eyhkr3o4fLwcYO4Bft39Bpx1hGnmR0xGN1prpwK
Moih/rqwTjDLBwms/rCl5JY5mJNIJCt6tzbzPNXOk0SXerLmafyGdXXm+qjDLMJtoJGvkLAFhIPL
PixDPtzcaVHf/HiSAoM6Mx6ekpBhErbOIpn/hdz9bPsTZt87C6RaBn5WULGsUsoYKYwGKSEDt2PJ
/BqflVzjenDSA7xv4GYfSiUA+Solhcd6btBwuVlDA7lFej4ZUp6LpL0K7UnkvcS2RVnkrAynofnJ
aqe7pyqTqQlM1NTxFp2Lvm5r9drKiC+jtp1+GIS8rBvLWcW2IulrOeHFDDO/pLV2RgettZ2CZyej
gjczBMg+DyzxLfBtgCsrxFKqM7OEmToIE2rjl41oltQNR+LQdmTLTSsULVf2mV0jkIRjw1xN1oo9
13ZpgVARREMzHPEpuoX6qTizG12+KoavmemzSjG2lly4PasvtRR80Py7buHjqidzqYOKooK9oiHs
g+ALnt2ninMm5MznU1E/HjB4oxJkY4zg7EoEy9Gk/pjVhpEohvuaXoeVYleSxjtpM3l/pZpWh4Z+
jj8/uHAdt7vnWdXyewJ2QSknn34PB1SQ2DoH7fgXVlOjkYjZpVs6HaXNHBoKYXEV51bzTuR4/mhF
ET/OIr2p2wRsKoGb3WEi8uwMePDa/b3lMSphj4GtaSL7hqF1JdPwHw/2eu96IchdbjrHFgoF8EPA
CbZD7kTmFA/afAXj8L7uyFZfE7gn9pxtce01UkE5M5C5eMwdpw3XYKcQNMrmbjS/2ZRvYZQLLoX2
X45u/6c2tzXGZgtGnLH48fIlU1y06PQXAPFFhkfQF1ME7NCF4mMpLyawZQU4SVFXTgE0DmJdLvuC
eafdpNZ1N4drBdzsCKsn5UNRGotZETd0o6jfcmXBZOlcrITVBHPZE0bLWNXEoo93nPpQsKTIDJlN
XBTkvK2KE+4Q1bfZiTcuj0JlWmuI3I+ZkWpFeLt3Pv1D8ujla2KTFEuPtWWGAtpPC3vvuybn5F8s
dNdicgqo38ZNV1gzdriZIdFb47vmGLYWTEC6xGwm/Nt9KwoOF/Kl6eegNswbaGU6jl0t2yBvhiPc
hov2xY2I1fjEN2KBng7TnnL0cQNMqN/IEPxg5mlMy0wE5/qmEG9Ql38UoH8ZHL6LVTPj3jpPBCKA
evpJOV7wBKdkCQb1voFn1F4T8A3Eftg8/6pPCz7k8C7spZgbgxuQdeh0GLxVdAn4G3PbCOkJeRXm
Doh+xz3z7E7LSS+5Fe+8JvB8uRv7ax+sfGJqsp9uT2mlr+UFNOWNywoeeROUw3oAUXpvFRrzaVkS
zKrKb49Lf6CGpFlNMzVKMMvAQacT2P5/Z+Ew9V5w8BB6+lztYAIHgXKyxhLjg4/iCP6MILx8X/f2
qgNr2w+Kh+0op609mnyLfewosSdcoiZaZPgElH7ct0OGrr5lekUA3e6ZLJwuVBZT88JInGnN4veJ
xfDIrzZWJn6IDbEvuuB4WYPsRdBU7mWA2wEdBw7CkzJruccFgyeYt2JvtPo4VwY8O6DYDQ2wz7vW
PVUyjZ5FeKbpczTrSbtTvY28KujINmLTCSyUbQfVZd2N4Uyz1C1A/24V+nzM2SOMv6FKZhbC+Fw0
+0qtcovbwCe3IrMk10/mOmQRMigx27JWslOlsEERsCRPDeQfaTql5YkozttzlH4zwhVZsysn3R2P
R6UzpdxUONb4hNSMzt5y7qa9S/U9dj1CRhd5GDyY2b9AYyPzXGqGVm/7Hf1KvaJpQJ4ObxtRDOVV
Y1J75qAKVJB0ruTX+rO+N0QehiHtEv8IjnwzTRQgL7xW+rL/1G1YmJPEZ3QaItCzpaUCyc1y938J
svx7y09QrCspJuZUw9cUFnOmodEbuSZf/GB7iejuRd26+/7Rg7oVNZieOaOywvp1rsDsPp5uHoFU
dvphdE/Gd9xseZUJa5kNPlJPad1KxOqyUQjkDQuQzcM/swZT8HSowgleOAfpaN+YutWQB2k6ZrWS
h8Kz6ChD1EiuhGuSz/b62I8Tann1YQDv6PM6THmsAKOCWhmEgidVusabYzACLx5CpThQUU8rMwb8
Jm+7BDNbAlFkq/53Tsrs5NqscNbNCMzCEZTw4SK7DuP+1n0FrMssubC1CV0/UfVCQs+h9BgYKpcS
PWfdv7EsImE1anVIO+SGwxH7izjiwUInaxAP4wbmiTp94Y7bTh60EpVy27tzXAOlLaTL35Sm/mh/
Iu7aLYpHUlQ0RBuxqR/XAgOZsE8cevsWkkzQIGtArFWoj2MI9z02z61B8K0qlXJXJrmgVE+l0ucU
CQNZok1wUFnTOHLYsPVEWnIH23du1bp1+bxqk7r7tiw/pQJxEqX0MWk9A1G2MihWGog0U/8leEf7
BmX0SnxjPryx5KMMrY7Rs/Xln+E/K4WsIaUvwVCdOkCHtjMJzRXvExvu5V8rcVS4d1aLQgOIuONr
ow/f++p7FnQ4yKC9OfFat5lyrXc2K5zy1UMko/eU4qb5ZVon96xr6iY106kCkpn+Zjr19MRNSCpa
ncMs3Ndvq/dnHBs7enV4fEcDvuOZehPebWyKX/XknIu9LHGQeY/mRCFhQYHMSn3Vck1cWxD46Zdy
3xShDx+/J4nw+EZVRpOzpHTObYvbxlVJgWrD7mneKjW+FMDtJmP8IaYG4vd77Y7q6tPny7Got2Fg
VUlj/zbwjkqkyJ3iz7oVNi6pBBv2JekVw6bsUnyXF2/DS63iKUqAEGOUnEAnnm/BGUo/+aQ1khRs
zJ0Oz/dxXCfDX9mtUCovzdF9q3cnr/ZxdpVlHFrN4UJIR7+wOvgdZIq9fQgdDknBuT3Bt3yU3vfV
ejQrxH323jNeOvaU/zRVP1C8hXnjI6oxRlkkXmaEV/qbDGemn9W13N4L7hkhNEyknQRQ+Po78lYR
IyzaejiS2d0zDouFQVXrwCUe1suW6VQg6uGmucrosGaKedx8hCqPZfTn6wy/fdoCm/mYtiVMfE/B
j+870mYkCvDdJsAz4dm31i2PgALP2sugdsWph96FX4ZD3axgtvJjJPbkiYV51sTOAmSBZb7v1Hhc
dQyNIDEE6COeLd7FVLe4wwxByIDLbQ6blgc6NawE1RlAmosB2EL8kilvWo0IfYYrzLDuIWGuTfSE
uX02RNa9cjwzzA+Y/n/jv57u8YtwRpE9EAqciJYIz6/s5I4xN1RQcfJqoFsp57XgjJzygyFeuI4s
O5cc8a2FMznBT4JnMkwc1o0QiCck5T/1CFWafSrtVIAiBko0fgl18ANvmqcyztgGRUomH2lu+sg9
2xLNTIIvCHX0FuWKq32cIi2+t38cP3Y06gPQtDjdfcGUMMR5Tqk0Dj1Ku748sIkrC3UDvdqRrQQg
731RCEojXD58zse8+9LPabMidiZqavnc9u3G//LbtfPKl0Z22AGRwMpgXheFcs6LFR/2k/d4zNED
JETZbLb7RVAFcur1/7lQJxaEKyH17YOnXXgvKPBB/6ODjmLTzEssi5QR4hgs1J8rdq63WlLx6OTN
MhIncF/mQYnPKS9/vvlIlNw457AlE0r85ojlO/hN3ljsogeMEx4I5U/b4d1ejJVtltNnPBw1YJZr
G4Zv8DhlGFUUypM420MhcTR5oOMrYu5nHni9WyAOS2iTHxbsI1QoYheJJUCeiqIrMgoYI6LMyHsP
H1s96cCDoeSs2bGF+GgUxvAzdqCkwxcrWccPMNV+XvLUxbsGHmH0ZtD9e9yJ8F15ghnhoPh0zpmk
cc1dnz4dpwVBkpcXtoVasUi1If80H/zj0XWYS07v1t/HfXioekEbUv/BMWOYgD+MT7LkHnVYwokm
tv+tALyofj/l3JLLTv5H8k+ddKaxdnHKGfbPm4pc5wOcudpmDbdWWsaZvYQf4MKwIL/J+wAU9DFa
W3qCHiPinZQw1wAzqoYpt70Avys3/KFVZBNOSKGuI4YFRzSSBlXMS05ef+xH+XXpCSgDgOftfuTj
aSW2u03u9ya0L5KxUvf6EtgL0pnJptNQZN7xnTHpCl20cJbP4D/uCAqys1QIgpAFS3EltOeKrWTe
qZtmJ5sBuFT+c726G4J6kOkpKYn9SyaUxolOKxJ4fnDznL/SQn2o8I7acioZVJZUwRzbGNJHEuB5
r7UtnzEkxv8wWAC2pMOr3sf9H8ZX6v457U6EWliG263EpDbI9U0xRB7ncXhdYwLAuudJu5Hhkngz
vA3X2+igeSGKDIpXj3O9EvVXo7pfLKSnYHUqoTrNrn3fCHqt6ykU1YrvKEQi0u/tdG5l/R+AXDYq
qqpSxHnd1obkENFrG9kFLdOSH8YTTANCbK2aQmy8RLNV8cNSVFPklHs2KUbBaHz4S7fBMROsoteq
pwVNgFgwJ9y9dVdmLIuYH78Oop1r5rvEQKdoHT4xpsrIHWIepmTwi69VdoiVmmjaY4vwgkHw+qAx
fHDG7qszzB/7M90bGuM+sdId+NrQ5j/2ejzt7g+PMMSUFQtjRKtplYv5ibXcrky2um3STFU89f/W
nbz1kRt4TpzD8FgnFIQ4mxW/iAr7YhlCvXnsR84QeMh1NW7m2Zr1I+r6fDM696ubqUEdU6wNvHxE
bjJXLbsbrLKJjtMTE/g9O9dlwOFPW2hEhah2uoF295EXUTmdXSakBJtrHvukYI63dJlgFkmhHcjg
6hkduV2fYvLOiW/ds4dM3tGlDtHKF2ggxIc39q2M9U8tY3b8cOVHYmrGs4300Or3Jh3+L5y9MZ6V
0iO0lW6C0rUhxD20mZxhCsSlmTkwp1GRtQCWEXygpjXZiQJMDSTyM3USb1NIfsyARu4qGBGSpveI
gZjrpH+3qmIEQ0d7Yv/8fof0cX9m16R8BeNYCyI+6RuPbc+MqKhzhDoTAkAWN5A4pjMrHwUaCGDv
Q+ZBS/aNjHYpP16rFlRge0PxVOLlDXqjGNKCqUQA7XN1EV3C+IKlI/+W4zMYzwPhfXWUCPtEw4m0
Ew2BDLiyEKp0X63YgayD481/vwHkqIJyCWOOsDEOgkV2iFq/Bb8HmyxpJkSlCNwnZPgcqHKRE0Ru
JYt+g+Evb1wjfIOLQ7z9yUuXOvclSwLRXq1Xnz/AHRD5P2wVKo9rr1KBR4PTVnHgKuiwpHhFVdnQ
1IxoLgbjW5mRCkX0fat8tdOKszNqhD8anS4Cbe446LrrgRK4y7qaZJfCVtDFg65vFzY01UY3lIdf
5gHk7/RjYTeILLZxgxe5jpdykJBywOCGWpXFt0b7cEigpNz6p9tXJLsJuy0f+vsFeN6Vyf+acfNi
MO31E2RZpXbK3puDJuonqCPZVqtgqt3clxNEGXJ0fQZvuNG0qSHVenYX/GiRPJnCTQDr/qVLvBcf
JPpTAzPI3YqgYaw/k9Lqr1SeBHqIOjjMTR2gB4tzmQXslf0xd/MzX65nGf1fSBnnzwuGFXLWGjJy
GmksuvUNpcBOald7ntV3ljPUbxyxNNz/ZHQ3YgsbqkBm7MMB7CjxoWdJRjUj0buL6JxqEuDofrwn
LTfc+YA/0TBBzi8ZfDXSqMkLavc+U+smiq+buCRCqkWfVE1GCDXF1FGX0NMZptlwF7gmmAI1yKfG
8R31ToX+x24breFMeSukQXF93wj7/riR7w8AiWFXmvErkevIxV91RdPu4bVoWQ1w6QDkcc92GKjP
YD+vN75NaAuldAriLHRnuHVBxOuF944H1GmGT0xo1y2L/ceTN+qA9GB+dcxSQnvB3vtB25pv2ivU
+aq6SG4SMuW0B/ZVaDi7Wb4CYYP9NHPXw4dJ3WzB90wS4BHMvMD4oE+6YSghRvCwRHt6Racpelzj
pSCkul8/GspPr9evTHxveiZ4CG0aEPUzBz8Kx77IbVX79ejjduz4+P78+HYlNoTxIocfriEGbBXS
PitC9QlD/BW6hKSUbaNiRCyDYAMsd9YxK+Dj44I8SNhW0tN+n5kpiYrGWy+6wv+4DHpk5v2P7w6w
ZKVAfa3H5FMgoqLmep69ofW9DCNYv1nDr3ABb4oZ46MIEsi14B+BoxdQV7UNO555zFBuqye4JqJT
eripHIOScktQww4rU6YCxMy5Sd7/59HrNYi0kxHarWyWQfuWVxRaSDx2+Gjf9WClhR73S4esvsx0
WV4ycp7k3sKPcmxgnPf/TzDjmkpYVsgh36V6OeOlfGCS5WGd3t1SO/4UxyEhesO6B/rtgJn7M/di
hGLgFFE9z8uylZHZ+X2PIFiMv7+hi9WeJvy/0vzbm5JRnMYfHG7ht3PWBSJK1jIdwyCgZleh2E17
Vt5oA8tI6FtTvUQQYyVINKFs1feeGAwj6oIHSSCeOb1oME2weRBeATa5qLWaGtMXaSyLgtu9fa8+
uoeM+3AHpPbtAzZPPfc6YJ33RBKrp7Ud/zZwwG+YgCSY3K+eLrRAyRIgeRM9Z6qrqW7z+QODw243
P4b3Uz8HV3If3ykNjb/dEP+TL9ZaXRwtyNpfkn7kppbiDR9eLQ/P4lwS7Y0GV5S8ahUIb4sFR2/V
Ghuynfi3rbq6e4+enwA89xsc7inc5bohdZN6q+e1grEHuwNLc48O0nHDCALPWXQy2jmG37ZlbwUL
YZ+JzCD2Cj97u5ttTyLkz3HUKV9rV6DoKpDVtojnfqF3sxE5OLoBPnxYZO8+MuYg1vqSFuyo99Yj
CA5mfZNekDVk20SvrEihE3s5FlyRA2/vMV3I8+vQZ6o9GV22HxxfbiY8d9Aj/dhJzSgL6t6RM0M0
mNK34z0OUsOtWYVo6nQsqvwjMOumICe3g6yZyYaITuFAR8TezPbi+tTugfUfVUHHb8z+H5rpUlTd
NFaLG8mwEwl8qLyjV9cwuRt1Dzwx+8S4Q7eFMS307BvMarEj76BPy6kVk75dc4uvkakX+2ySy1la
UVwPRbLjQZdJtaBWabZPYhMtsvwWO51jV+ua6N4lWNc+6Jvo8GhlLcjVVe4mFWKzVIH4dVro4qZV
Bm700R2tOHW9wZCkYSJoL11bETg6wxCg+k2ZTMSo4AAJcES/Tt5tnYCzfnO/s6/54KeuFmVOZ1/4
fVYN2kGhnS4V3Tc2Lf+piKjqHIiM4Zxv4fj/IqgecxAUgkLTgpttjAcTiM8PTLtQUYvssSpXR4am
rQalyvhFHiZGzagFmI6klxErwRmZEOvWucTXevFL62OKJhlOQCSBoyb/1sSD24GDrRYkf8IJ8Nwo
9Q/riJ9Xx3hVWI4oYbAG2Eavjl/ebaNxxv3RDu5N7yLyp1SbBsvHtHQp6rQBLv3r/MYxneFGJCPV
SqC75ttPdNwRyzW3zOgDEtyzsxbuv0e26pzW/8b3DiQv4pwBsvfnx0YnvoMzBD/rcezczcVbkhWV
jCmHL5u7oxlHFuLlQmw/WhepkgCdDnzFjSQSykHxIiSIQl+pfSoPAssgQYAmmBTLKUBfPIrt4ZUo
hJ1sCWwiWvsQXb5/+Qnw1xnZNCFrISdQ94ffS0pM1GB8Vy7PM8npl352fG9dsda2iDFWT8ezLMoO
2nNzSHBiavZExRZNdXSl9SyJdtL0k6u923BmYm2r3fsOpdW3Yl0Os9rjWU7pqp2hKgNhuBZKVUQ2
tPSIYDg7+OzX5lZZ1CzrNU4zGKwmTM+xpdF+y8kAjvfCMyOEaU9AZvzTCeEE0zP77dNsTafJI5pS
Adx/C4abCyUtXHC7IqzBvfgf8m9H4Mna1RDwBy1rk6XaD8voscoMiV5vfy8L46Hc+i1B+i1L4XF5
TUKtYIC+lFIPRRN7VyiQo+R9KIf6nMC02qBDBlmyY+BeLFB1bs2RYqK4biNhlA0c4+BYc35hChQw
/uTVKop0AMHIpTqdkItzRRUkANaanfZVaOg2x4IbJUVZXxoJxbwav6phmlUKkrTeXrY8ejyCy5s9
VSKybK4ZLh3BawBKdc14hjbnJuCR5idCxbHVRNVuhhCM8gfq9Tp/F05eoNIzO5RczGEuWcZgI+uO
s+ZAvDfqoslm9uD75j82pzvg461mctpTavW02e4ZgtGhCcmOm0bRqAD+2F7QgFa10Eq2pVDOUC2P
+vMU/ccdc6QTCI+wSVdvyFrMgxILRqyyCJFvtgvDaH5HMuElf52PCQ/Yvwk12q9qRdH20HVXodAh
hw543VO/D7Q/2vrjM0gXIx+2a6wyBJtQQHo0JHtffVuyUbzPpRJY25dT3WkMqbo83rLJARs1GlEr
LhOqidi6OQGMBrEgyx1qtwAhH8Su4+YNpiYPP8P5fGz3S0T5Edo60hhehT76Z/AfFuCZ44KTZQn2
lTxUIHX0hFbBTEsuzvY1fgm3JrecvcKjYJZ4VR4jCxa36dafGwvCwNqa9wg8TCJpLpCJiRGFW082
OkSHrxE+tHmpB5N7PIXrQI/FjpKLG8E80BPj4ZSF6I1S25O3YapEVI9Txru7SAiMbsp2yAD5545s
//7olH+GyutlXenAX4LlRB8Shey8hmJ73eENBKnKWpAADhAWp5fubk/NIcD4zrNJZkP/g9VqNdjW
67osNnKdbu4P1CNTYAn/7euutx2MCwsfSDC8PxX9uNWJ2VfjkZS/rSpm9s2M1pO6sc7PYHtoRpwe
0+5tZYGBp1XQLyZ5rlJwbkyecnjFsUDZAn6gzSvIpmAG0g5Bapy7HniACb20Z8/xcLPH+YeOPHgV
2HC3eBFRh3rQowLbWw5R4xywVzF39HPwqvkRZprWiE2hR1Xm6bdG9ICVXTLLAHbJf9dL2oSGEd8f
lVR5XqTu3Ix8VfO6a6kaijDucBKyPAhUMJDvCDC87C1Dt2ML5kMGQ9E5nJE8YZGHhks5PVkvp3jY
h2TWSRabMDdTpIa4U3ilewU6cWXJNyhA7fM+BnBzc9pn0OGa/pnYF/oRR2alfJzR3tyRWLW/WmHi
GkC3qJemJ0XZ+Cv7R3hzFC6st6uaKj3kE0mDC3oGephlNBZa1ZZagxegsbqXRi5NTBwnGOIv5HX6
kYTTVS7/ggBPSENR1IQZm272aV4HEtGCiWVz3ziNFiu4znG/QWz44M2X2a/R5FqFhm7iGsoqgFNt
vyLeJvPc9Ie2CIrO64ppZ/lk4m7ojMFwGaC4MTs7MtoS5CF0mp7LbD16Fe/+TxGuUEvm5WCG8BQT
7cJZ+Rs/vCLjz2nNL2KZEDxJyOhj2c00OiklOu3C2ZckQSL2vFuC0FUgFoTZg63nT9nEnDbXiPd7
8vpN3jr/rVgeJI0zzVYd144yrBb5B3o1hel+fOt22eBycuMdil5qFe/KDqaO7FOCuCWOPa67XJor
DPgIukiZHhOdEXEkFaKgXpp4k+3NKlvt4cE6t7qPf0JeuJYVJscabk3Hxrr67MD9hrErzrRbw3Uq
CKCjytqQn29X2dsLIrZtbcNo1wfMPEHcRb5aqwS7hE5Y7UUqMvjLzTwOSS2Pq3FvtZCSeHsNXhmy
otC/je4hSrw8j1ngadJMZuXurXo5jsB3Nwg4XWiecifK2HrG0aG4FAcy8GN2xHuCE+Ex8PVWnrGC
/Q11IDpw+1cySF6UEn2UCh/JKapRRnIUqPSdwPDQzkgydl9mSonejf1sqhiNiic9Rd9YfSbUPeuQ
7H7X06R2SpbgXI+pig3eouVM4nvtv2keEvDJaxuIblqHGS4q1x726fLeGrHOF+hNIFqUIuUo9HCn
LL2Z02LfCqc8WsWd8XO8CMcYblBvrJPpVfaqfoKa0sToMX1ZQ65LEscZkQgf11tpcKGzVjn6ynFZ
7ccqbR02t2FrdKyHBvk/oidgzX0P+q0TqZnwbGDWTSwQgkpmpMlK/QycCX/N176z3x1TiWBI347l
7ps4DptAGxxYECUdiHbFdnyf589uQSfckfcj6ML1OSKWcJHqusiyorMRVbkuRqwhiKwUpIdNOi8Q
vxn6YRvgMmYgSzDQzyAfxfMMCPjcVlf5ejXUDmLoI2yr5u54l0/StkI2Xmj/NdadINRFtao1Z3Ld
yS3rWueNWZavxSdMIyBCTfMnSW7+XWETqMYhYcDZ5cRdC1Eo/ZN/TuPPNeCrhgMDyZKK4Tev0Oxi
yWHgIucFyMWXSz805o7KIPXdeMb5u6p6/2qCQMsvQASv3uZwCux7pmf1h/HjezlY9pM005QPZDEh
kZiYzUeZnssrABb5RA5k5WGA58rNEbniEZ4fCOHpFvd8byBPrRlzIk5EgJ30QDpidGpTmCStAPO/
9fKm0z1+QW8VeC1C3hTttReoFbdkvJBG7k4Mc9wFp5ebD3DAtpBul9wzl/qf45AxZ3S7lCgOlZDY
9CdtQgjqWkTAP7xsTFGkUF2rOfBp5ljiVHUOVEdOhVBjWzuImKVoUhGv7e74lYjLoQWpklpDbFt9
Lfhgc+X9lQDlg7rsIoOOCIaIJeWJDuJKCdn1UcziNmVhwyuBnCQfIJZjXkc9ovhqtGvR6HoYXrFx
AIEi/sk6LhlC0XOBMtU+ORWi54xs7dZG5tTGmfp+3PYWBprfHmVRzeE0eIQ4TD12cEVxULwafTyR
hj7lJ8M1R5U6De6TfxcwqoDbjyMNQTz9g9Ios/gZB0wuX/X1kILxP+8JGiCIOyqQJcpzhr8MazVD
GqK+piGJbDrA0CVHqu559p4xY/ulLK9oWO5ZrHHrOz3j0YQqCrTIkKh5oqODDiDmwIHiduN9pt3L
ybJS5ZeHj/6KL4tx1BK4aRpokC7K7H2QYPfGYt22wJH+e7DRcH9g0HEuhmQlM2rBzUiVHYCXaNpu
MXmj8Jf2LE5jMdJE8DeAPy6BAa4sNpNLwhPqT889HEGYuCMyewA80A5ji4QNWUkXIAeDNQ0lFUOz
O9XdetOR7wEYs097XKl5oub7kdAJe23KTzIt7E4gPZ3XRAw084tNg/u6GVBsSrzVrqCLbj9h5OWH
4R7exF6VjE8NsOKfGpX9Jr/I/Oe0x85Pyz3Kgf+ca2btNQlANLqvMtjHuGgQ5xU3fogANki3YIG0
0sI+qgGplhXrvK+/2QEKL3/3yLd5bvW14BIU0/xlYzLFQE4FjgVxbYkULoTffPgVwDkrE8PWo8r0
tNxwj58SHNJBsgpOShjyxPCHfruIoVJ4dNPWWOTJdjsrNmZGg1zMD1r9W0y56Q6QP1q+Rb3mVXA+
XrgnPUuSBM3UBqpO1HrSc2+kVVh9VmOHQ5NqSNJc+8LKtex72fJXQWsrGdotMpj0C3OV4dOrqJ0l
8OF3M1h0fq2Sgyds3sc2J2DwhYUFNN6yGytMVJrenSYym2oy0XkksgHsTlDewrjNAQAZ/t1fxd3H
JBRWBez9PEoGNhykiTyaSUwlULR52mmt6WJqAK1XbxP/+SrzDbGR5X/UxlZORSIkSdBnav1IMrkP
81hcyObonwTyseoEqvKiuGtfAvIr8+3M7hAVEyvCIcQ9YrVmn8Tupgap2q0Dlw7ukIt9uytQF9f4
qcgg5FyiHxY5da7htkv1AYSRTrC7VLLfawEUwsuIxAEfzRBkDYI9MNfat4qR+6AqabVZp+k8O5z8
ZLXnIgsMDph2qQri/2JfWCcwQHQUCmiX+GbOExHJnrDWzQ/RHifQfx+W5VTEFAVLF/iKaqjKZrTB
ykIzekIqx+SXAHOD8yWWvBbBXnTDZB3Ni379V35Vt6ByazZYRJmMxNH5nulKykWQYbg+orJH93Yo
3LZHQ7BGTnEd2cTmt6YjigcqtbzhU5/Y50md8a2EG3KtHnnaRRa+ADCcRN2dXAwbSpqNcd60EeyO
6gzrfblAwmXILf3sHQml6GxjztDQFEix4uyGRxoMiLbKOYsUooGQOTvWrAzcfsbjsuqW7ZcQDOoq
N/nlgkZ9M0u3LH3rtOGhvfUGIujgNgo7mFiJB99xTylc1vCl8J/58TTqPa4SNQ4tr0Jgen1xbZhA
xZBkH8XxFjG56b6ylQlWcYsNRUNP2fMq30xHtz0akH4JQ4nekQTEJLht6oInOJXzDVrTSqOrg2t/
rT99x8ba7YH0TeeK2brfUwzU3yb4DomhEHuLtvcb6d4m0yy6cKAndHo+5Tjt2KEIEo6RcK1rAwhj
vCEeLRCRv1V0sPkni/B/vJByMhhGvq+8/Rb/23MkfuBUTJT+ApBBwjnod3Oxx3huZPS721qVmf8X
4gqBOnYjkNVfAMBtzFbl4g3CjgO3dtw5yEIO0LacM68d7pu1wv/25QQBt+yWh3DM3lLdqLS3tjZq
6QlB1kmgvXHjYd2fLacdDZzvR6SOzwo7uQUVJgWBNvuiEYnfzLYAwAej+Ey29rHNQYEf5GHQss9z
CSu8EgjVU3Cs183JL/9KNQ9VNQQSu/xvu8g136iHa/4TVOsYO3WICiksEqc4ZQgMAqL8B359i8Mp
lMDisgakn+1u2ia/P6nXWF3//FqTZNp/YTa61XBw219XQNybQ0/Gedo1V0BCXwGPURYzHbnqb5Ks
3XI1piXQrlBQQuLbqZgv9r+Jr/H3NlFIP1YaXCqrh9Yu1T21nYtU5xv7Sp0HyD7sUQDHj/di+4+q
wuyaRoeWhPg0M+MbQIc50KAhSFRCgMhAtc1Gn5LOY4RhS2ZiHuKsQtsedfytLC6jrA7/ObCbqKYj
kh69/0eNrvmU9wkWLYP4Tv9DDjZIuF3fD7TyHUTqQ3wXaThjqkSN8EY7s72GKPDYIwM3rvBmh4Ya
1dDQFss52mBliLu3tAM5+nBzLnjUuZHr7OTHkksFd+ldZfVmfCZIhVdJ3mcXNQxBXBBnsZdKnd3i
JNpxERu/vSdZTzHY+GL8yIw4yIlvCIRnYu6sarrn3yEnpNmxNVaxAoAVtUWVgciq9E+34jWJyg7h
hugjRd8mSSOYAKcr7hwpuSg9CBnQuMNYKNOgcB+/KRkSJbRKqC0htIH66IV/KjnIMyf6J9v5HDlZ
1ndzJO04MARUiTgtY/cGF5F+xXmSZiRyyXYi5XgH4+HB4UzGN1Er48xF4utdq7URtCP4YPHXuOqG
8xIdh6Ep+yOXINKzrFjAOVZhMNZcQ4Y38eD4iVB1CyxPXdiKeiMuAVrGAJ+gnvElM5f09ca2hQ3c
DYdRNb+SrNucCMVBsqcT8b6OnYcwzFy4nXIKfwldsQdDos0+DwkjTeIJUmjfioE/AZPikxQEioUR
CiXgnJiyAMmc2NJofkwNqirhPo4Xyk4/xE2sRZJqwSkpFB99pGN6Tm5s57DhkijV9IupraB6msZw
IhXZeQCTrgeVHNmXoVmOe8kVc/MFAywU8uPLC/bRV3OkiwHiCufcIAdlabBqltNB79aQfUZnzsUr
q1Spb8nrUop3VIwx0AWi074BF532xF/C+uE0xnLIDf7jIY8ryAKcNpsDHck57MFT6xVIvJs7ImxX
CtdtS2hfzBQBrxXXEKE39C2CTS0iNjhneVesXzFMVd/PQ++BvooyaLpieIoqbFe48VAZPBFkiljQ
yIGR6GIcetBE0QfhJwodGYsEHCE0DbNHYqqcxPi7U3O7ZSWYy7MsIJmyIDYUWV62gH0yyql1U8+c
ZUlAkZK8Q6tkO4Xt3lztm8w5EyaroWWs369e8V8KdXOO8Oeqi0M1vEqmqtZopwKR1gB50qE+XN2h
gMru3YpfXOVUHOT0W3H8+ILy2u2ZUywt+33J6SrtObLPoALNg7WtplA1U7zqmUMLcD9lepp43PkM
/YTRBrMY33v6kGklLF2+E264F+YnSbI0cZbyGQpikvSgAbf7lecP6kSnYhjDOmo7eFJB940X7uL0
eQBOvIl9lrDtoy6nZux8WHJ263KJbJPlGrufvJb71lPLdew7BSu4Ln6dzSuhgS84gezpfKQ8vofo
jDZj2nobJQzrWwNsOOWLvmkaa03GGgTzl++UhouDGUjoU+6VMaD8V7sEsHpOUj3aRe2TSooHl2mV
GxyIbyOL67eBsge955Eph6F95Po5hn1LHTN2foHPXVKfrhipDujhWcV9GB9CM9Hz2adCzPdGm8Ig
xg+gG46qK7Kjh2Zd3vJJZEsO752jsRN74Ud30SuR+zyfDikGfuLgMsGeydzXSckvwOIn5iyPD6Vd
oi/tnf5qhmbmTnYmsR5q2WIx6KE8hXUQXo7QISCh+YqSdfATDMIDtilE3oXy9/LMV4jFlaeOWAjq
hUyhuyfyOn5Z5DLr9HNf0TFBOtNKFd2NEv0bCJzn7YqEhILA8qKqAZ69wwxWN65F4uj0h64Uf24s
3WvQBQbc/eS9vnJx+Cd8M0C6qwOZccNkF+4i3p/4KNDgWzik4XCvubdJnsNymfjDukPHKY/+IJTp
ZrYyabuX5XMh1a9InFD3UydjLd5XrQZy/ocscsSUtOWBwxwgXHJwoAzzOvbRHkIgS9oQtBphMjeF
toBTA0ak8qk+8HQcZDmcTfaERH715ZC9P4krJJbFkJ7xGxQpMxokW3Pxw1/IMDIzgkUh1Q0ttubS
BMB8hQK7cLtz/RzAVwpyMPAcQ1B78+YOQG92LKNzO+U4PJLk8APavTws/qM3x1Vio3S5Pk4LG3un
8l0CjuNirapOoPJahTw2fBhrNkE8GhmXl3XZyWKXNlj7Z8wSmTbYtmlys7sJfK1tUqucjplLAhsg
d733dZqMMymTBgon7zI7V/VBflSIlA6fyoKJV3el0P2cJUHd6p3EawZfBy+9lWv7LY7sk4piRbj3
I2RORmz/07BrgbsLYRkfFO7IpsXxDp8FFMubo9WZ1FKw2U6kdu9LMQGRn+amPLx5xUMzQ0d+N9+t
B5msuCJVrz46ri21kq+1xsuzUCcsXmOCLRW1IfmtLd+MtKiz7wn5uiTwSYIRRkkAMsB5xtJ/3I4C
pW7CcKC2H5smz+1RhbWm+xNZqpc+1EjxguYM1U7hfnLRQH4PLMIgYPiXaCanvF2sV+Sq6Q+nC4EX
DqakGYH9Z1rx7dEtKGRi80qM1htFM7zuphd4PfKP3ZyQfKLmH2qwiR01iv0553sWSW1+u5TyBMP+
EHbeUfdwKM3EjQP9oUaRbMNv5drugbrBPmJb0vSdF9SZFFmVAseelpvGrGG9zwYylF0IWAbe18eh
fyCbO3HaPr6QrqH/5XqdesbsniO1EL6vQOiTZnByiI7eT2ShyO3ozyMtPohy5xuQH0l69bjWCJuQ
4oR/X/mSPcG/ybepg7l5JRljPsp0izbnD6Os3hJUmwLzda7ow5Sg9Cjj2GebQKN1aJKvhXq8hqjQ
GtP4dbpyf9P0EZQQzLxSbIpS4qLKy+2UDfgV7gGGKcjq8tkbWrdRtqnFxHTUIAOzOqpwI+dRJB2e
LI2YY2GOd8VlCVn6oR8iQQDVbTXKF5rrnLvdRoqHmfNhipginc8zyTb9BD9sESmYiyooPfnIM/7m
ykq2jNHypjHy+DE353/YM840qnWaN2heHzTlfmoMS14siLrG6fSuZJmI9wF1SVLAEmqnb8eWiU5+
An36SceiOrhzv2DYXwzrPhb9hPmBTdZVDA2WHWuoLMOLah9vlYRVp5tIV3I5AfIOgqIfhDucqU04
gOXUQLZZry3jeyKLBdpXCXacFqyAI8O51ZN3hAlFqeI6zfbA1kuw4iA2+Zl8BVLytkExzlWxlBPR
Rvqey7owTeRIPfSgNdFe/rX7vGryiFkRj25F0L6uqNqanb2RtPvL7aGQ+ckbCFETlSf7aPOAzjLK
Qhv5ZejvnLVsX0PaEPQp4iWdj89ur+FBSb9mSIihp6zplHau133G8NSLlT2U93q7+3QgEHsB52Jo
uVX3qZTNRK0zH4Ogsx15c/g+FBfIgPz7gpTkTU+yC3h1/yJ9ZDSmxNz8Eu5mFg5XxOIJg5iUr4FG
i1WwdVbMu2JpesB0bl1W5VAdg2a/J8MOqIyIFtHmdHlxraU6G/l9LKhA13zd5E2Tv05xKK994owL
JA6YEUxdEt5a53BruMftFF3CRkb+plBQ099ea8K7Le7IOgGQehV+9kWpcsTay//I4i6gHr+aiLKz
tqqX38qBuabp0zGo92Ntyh+rQbgNWHEEV2tEEhejtFgEJsA+YwK0ClDjpPVXud7Rigne+m6mOfxJ
Y3j3BCoh7kfsLXY2PPDN2eVaYAGfkbhIaDQMni9B0iQ/owypQwM0DwK1hrZ2eOKDk71SyfK66VgI
Xafc6cRNndpIAfy08ZY294yFlzK5DMlOqQhTZ58JGRswLh4vrSPFjEe45u3iMvKYTOyBJoODiQw2
6AZrSI8Esdnbo1Din3LMReximVK7yWDtYvBxFJKCqDE34apGRus4FM00kVikvb2AbrSEWL/BYsES
E4Elkrqy50QvcgTxzC3olocSowlKJWuxltu80USvDfY4pKa2qoWWtp5RYmqb5cQypdAlcU5VKQBt
zhiwz33jv5dkS9STGtUn9MvJsZBMhUHpOA5jtu8P/+su896xayMygEXm+wvnfn1XbKR5Y9f8nl2+
75na+6gNubCLU4BiP2xB1+gHK2W0g+XbV1yMtU9exB22F9yrlRGvTjkvq1JRxXwHhMUYVWMVmymJ
RQstv6pqAlo2FTyXkZvUOTbxUtisFN3t9cDX/On30l8HqS2KhliSW7CEK3Qo6MJMz4+jdpZkfWpq
rjpGBEj0Vs4Jhem+EPCZGCCLe6+8pc1vkM45NAU10J8ahSD2ruQlAQLwqdNph6weoqNIk4QYSnae
HMbt7klelNlojzLCQ08ODMZ18m0egWqXHyvDMXKCxXFpycEuq+JQvJRcKYukFr/XbJfp/+xc/Xfn
yDjRDvN1DfZFY2wI0ZxwjofzBoqAL4uvAPrVBkP57gYKrsUA5PvTQK1W0YwsRTwX7wZiStcWxGDr
G6Dz4WwvGr4ONf0NdjpBYzPPL3yAr1Y/w73lTIKxnsGxCz3Ij3eOEPx4+ba1OHHLxibg7nogEul+
zA+cGCI/NTJA5fI9mmhK0NhOvxXZ85mxWVyYV5Y4MRk+eaubZPkYSF9YtTqx2kBbsAg9cdSUM1x3
MaF3j2QhjWNWcB6mKqAZpHOUbaU0TQ7ghCjBnZd1kmtN0XJJYfEguHwKxSUUaFsOYS8S1q6vH/aE
wo8kMK1LqOMAFzzmWaySE9I61PMDfCWYtVAWuRxw4+QEep6mYjqXeocVZSndSFcQcqdQ3vG/xbfT
M0ZFHYA3ph1Le2+mEw/Ci68EBymtzWCrnWhfl8spgJPNKmIWZv7wOiv/UXRQDXaZJYuHKTpWqAwP
1g1tF8H1NJjcKCHUAWPS2h+mt+9ilW3isatNPLpNCnicACRWQuw2qs6mQaCKKD8NVizP3dc5yPxw
Q6F4qx/GRlN3/+UHctPfQGONgTfVwomTt/P+TtQ3CvPNVf64vFAZs2efLBEmkczAwltMBU+5K/on
wmPNldo3jf4jcw8UkXt3F19EUuFV2HeCxnFigP08iMevdiTyGKWWDITcmvEMuyXKGy4G4ueLkci6
/Cvhhz6EBtqyMa78ktH2V3TKLoS926KbwkpiaVeNMX4goRyqx+SEjbXao2da7g9snkzIYXYrhGNW
vjtm4mLunugXx1bUo2sqsaTsAtLvgAIUYufs1dwdtqQzeizJxuKD8db4mVdRP1W5VkK1AhTwrWsW
Iag7MNkx6YcBCCzHd4KfryresWnxsoWL2J/Tf+kAfxwJu8EYCyOfqfRvm0o/qJjHM3q9OVItZnM/
ajdUMWS57mNsKxOIOoNW1pWnmYqutLDLeiQ5+/XATmrZ4L2dUAl4VFuACq9h6ESQlL0mG2xmNaSs
ay91HEjseZSkwfxqzDZjI92+d4M/kwJop1WEPp3zWeZJM6Yn95RGK/jGZmP3a02hTi4IZhe4GkQm
0iBF7MmPYMYOUlXxofclsA9/VCwxZWlieEHXVd2I9aPWjfFq52yhHE+vdBFiln2gFR7WCULfj6ld
LvmsjISeLl9EI/d0WEEHIvkjEW+lqqamsg2rdRiAt0Y98SYGAx4LeGAI2cs0epa7a0dC0kbuEVRP
UhDFPaef1oXuEqivqtjrdDMVqRN8jfsLUoUmclIfz1zzdk95VYL4hS4mNA2dbaRTM1qU101ECU94
/ytBJmnwFv0FtgxSIekK263KgM1cxAHFNoDRjVc09xkZm44DWMjQzYk6herBD506PlhftiAmF3Bt
0xmldcvzU0lYJL5oLfyRjMazx36fKdCKKKLNL6X43g8jCKBnXK9NC/I2A10kN44wmxNOdQLaIJSj
9ccO38041jpcxGW+Y5ncEgAS51ShKMi9H5NgXXC7TF4BIvjXmyYmzaDMthRm96Aduj+cCThT8cbs
i48zUhQFLWekX3/5NRgli9nrCkH9cCjsEq4huPGSkDJPAOiMAaQKiTCAq5+6tjvFxcxEZOdqrIVV
7VjAUgsWQBJVcIGFuKeKF77oNUjHv/Cz85yALxLJE2S8KxK6qHvxhb62vC5R3hPbHDbzlesrXZyv
sjMk8LfDYfpx7inCgMlnBQINErAv0Suem5akRkna4nGyPmS4zRDewljFK0R80eKmiFQWEZXyiJ4a
QUhka/Mqb0GFB3L7hmV2YFv+GRts2oeAi7ZViBuEiVV1t6HqWRBYDdJK9vwCW6AGm7D2BTLIOWak
NBn1hlIZ2Au1af0wDLOeSu3vCekAl5iw4z5HVgzh1qOz7t6mODhh2kVvpgSA1mcxwpb1TODV+e1b
JPZpPNpgP9QbjVFZ3lD/dJMux053NFdW8Qg000IWcYEe8QivIGecIXJy+eXWnjVdGokjqB/GeWV7
2xhVwnSV3c6DutNM5qSDBvRqSJIF6FG3RoH88R0aimJctzqnupaDs9M78ImLrulubYDDNlvjkGOi
+LY3Vx7P+6igWLtuZZfC1n6wAXqdhwN+mtWhHqDNW9duxG50w8KD8CmADqjkxXP7zmEwW33tG8jE
xeF41m4Tlu2hu9Qdn8jtPkLC4roMtFFlLHc0OvpRfgHqluLwDDBcxFhYxbEEKQR5GZolEVo6MXrh
89lW6FqAjx5nZU9g6TD66Mqb/3w1ahnhFjphx2HPkgD+dwB1EGH/L7cKOGwvrslP2nWGF5ZM1CYE
AIG9i2ASr7EbmDrPWu6LN0Q7BLd0YYfHXZWk52dq9x0ZK+mUPNRWVv0B+OR4RnCuIboh7ZhRaSCO
zONkj2nqZ/OaJhGLoiUmlMh3WiNqrdhpTCKT66icC/gkNPVbJWj/MfkYptF3intbGlNQDpvE99lw
AxZcf0IbnxcNPqjxNEmCv138IEKWn2ArScCNpWM6czgTTNUQjs0+7MD91xih8yhyzvZsFHUcGbuE
LbmmeIw1MTf5Fsd13w/o/IXxPwMn0FaKo7NpkdK2A4KmtzVUw7Wj4puWjXY8aUN0v0I6xvJHKp9p
FnN4VCqqoh99aCj66bq1m5xmFtw6049pclh5nTgUXt5kA3k5anWyPGG41DJbqMPkwwByJl+HlTOP
nRAmaQqjnre0TUXkZ2fNeR257cVMyPvf94DrrXypR2ged7+oMF7WhH3duENbnvM6PWKgDjFScLWi
LVBJJE4p+hqNx4BkVGkLHimlXRuQ6e5ia+EQ+XlvPSauvC2ZmCjGr6YsP14XKP55wt+skz16ejVO
kbQyZwncabCch8oLdb5dzvDHEAuufpSuqwuvgqjtvhpZDUxM70jSgTV9L7GeqlS3He8p1iB+HjjP
KYEnBWSaNFoZrE3YGwNfGhbRubrauEJXrGbzZ7A1RsNiiRM+1IQMeI7tMLkgzQg3h719yVNUAYo6
gVNgYLrM6nZrvZTKsQxTVq4ppub4acrAfl4tEMHZKvAUD2QUQD7Fc/FtXJEfs7n/TZQIrOnr32Pt
arHlqsskZIQOVBt0nqUrgO3tdwYP3HcBvTIChOyMpPar6ah+CjJxLAWHx4ew6mSgwsy9eMA4+bxf
IIdQIyR09AAp9VN3uEVbbKzon9DLP9XRE8JZxOqKSQJgWlziN2Lv5F61X/dPaki42zPfwT3pFILj
6Fl2UVRU4dMV/PJuMmtslChxS0KVYyIWD59Ggt6dtSHpR5jq5U69eUPgbdMJ0tUhaprXK9+6BisV
NbWasBHhdW/rr1wDsTJ2kldhFProoSnPB38vSLQstX07Rf0aWQLSH6UIn7OPY0U/+sgwy1RNlt09
PyR9GayjRrCDIOhsZJX3Q1Mi4xUoex6N2Ot4+t7OEfXxv+GgROybY3zROFqwz29THpkm+ypGpNlW
nb1iI8Ir0BbwgWCwhGbfx5auAoD+Dr+54cOR9rMQgw2hpQfkWKTV4NTWmmKWPFOvL9ajHZsfoDwY
Rrqb44IFmINe80EW/zVielhWNyPIQMajr7T5RN8D+hmOE9Lr3uFrlqZVZH16VlgTkyk42tkWe+jc
3efAUnEcDqkiVmkLbZ+M8FXj0KMHqR8h2HTbWXWZGlXh/oy1OwarVTql/6L2260LYzNYHIhMvoL0
9pQDbrPBMbOYZfLLAznnxU6rcO794lCjnqh0kIDwRv4+1ArQN7hXkF/oHLPjy5L9GBvJxrfXUwId
R6gRiyocKIjxq1oCjjm7D5SYPqgxzLOtjRe165aYLL+N7zFxVE9Or7HVNOoUww2h07cfN9YZCe+N
MTzQFdZr2eI/bWHe5koC6wS86FKgeOpy+sbkhxVB+3QnmwtcnSEhRyaJ/63qyctJsTeJ+lpf4ZdD
+iUNtcsY1QDubzvN/UGqfPkXtdJ6AKZUqsLb3pbnC5QxOObXvkMWz4Eey9bDPfNYSiOaRCXwFONi
AV4CO5oITfG/8ijAyX9S4gfGgWRGTrP8XxyOCkQknW+MLVxMbTBE2B3fjSX23Nl1g07Ff7J19Yhh
PDgSJl+1MTWt33QKxg1YiznZIB5g1sqH4p6bhIpLfCoQac9ZgGJ8NHtneV/YQq/9kBUpS11ZFntW
pRm8rYE6KV93kz4lILgE6qX0yL+8Ir9SI/3koCDEpQh7ovcrr3xH1A4Lzf9dwsb4+wFD8UoB9yw6
dPLCuHT7IWAlBFt00m1/Qctx2yGY5zBJ9rbVDVIEOS6fhX2mTpXYu1/4S9i//kmqK0vT6zHYwQFm
ij887f94XB6lMa+tt3i0emMYWLUNL+oHGAZX7ZgVEzpCDaP88VTGVcVFwlQx15BWH9JhdHIaWnG5
YEgw06wZG9nSYZgD1bwpt+J+qu5XQqxzj+p7ueO9gLRLEb7F7ISurp9KFLgY1uFd4hapCquEs8iH
CNGeGG3AmD5nF9c5vU7HotKwYUsRKOB3k+S4HkkzcISEZJxI3lBNPIrE7+DlJZE7jkxjzyFAop2v
L3QbVpX/NtdkpG8zpl2Jzo5BXFVW5EOxVJawMJBqMGHX2LZ7GbvDi/hgSJamZ+2JnbtghgJNc5lV
o5XAYGZ0OessMs00f09bDg114JOyDv020FItMt1q2IlyH68APOMDWqCOiiiLQfmtTBF36LdnZ91D
RfIpVtozgzxG3/I3pm7tz4tNb3GnNigEYfS7oCwv+Psifjo2STBTH2GE1CxzfNQgCHpKbMykRJ0o
8sa83KyMeS7aER2kSRA1OdflXwH5Z1D9XMmC5D9Ti/4v88oUM+MEo2+lxVJ7ZQSgQPBGv3IysIhk
OQN5ESdYkjL/OX49ahWtl0ioHDYl0rnnk7kvtZ9hIVU+SXOAAAQE563JuHphLWej5km8ErTuJynN
dIhR9/GGo/xbmSAEm9geIJ2s2EYrU3LQdV0FBWMqRYw9KNDKW4wQJnPDevLohXSWeN3LwcAOEwVb
Hiaghw0qwmsvGf5KENgw1tnH+nsuf+uiS8/Gta2JwNGpnlQbibs/pyNLIPaiJva8SkoPzJ0dVohT
tyDBRNJrenwYPT4i7KGTIPDGL2uLQt0bg0s1fHQe334F7SxlA8P6XH82Y1ROCmjqdDMbI1s8XVpn
LbWelJRZGhXLBQNTv04Eto+bmuHyR5swKYaCYd6kB3eVhSJyZAs6BWY3L5vKug1UVtK2eQ3Rl1eq
zhcLqmeLLmSdOfJBRGw0ELfAZKm+cuNT8NmFZqO/0au7f7I4HS+sFit28WAWlQ7717rKCy839Lzx
H1809rSZlM+6yzJT9Nf5JrV6a3Ayhxa/3L60xsln6zAzeNGxKqsIjxT8xGl/wWjQ6pZwWAwmSeLj
8K/1d2kD3iNvDrNgPVJkYFvIcOWqycaKpy6KcmneeAQbPdJF6iAh3IOPe4K2rJvcwcXSSOd0QHz1
n3jgS61iWT/C4RZtP0lOILKlEnNJ/CQ5LdutybjFX0vedUH8d3/HUg9W/jbN7nnH0xmoox7tEkR+
zhgWGxloMAWywyz0BFcgQ4dYXymDNz27tpmMndhRHhyfNtsC7JcYjDY84QHkqZP0dv+7+iw4TbtM
N//gFlj9/cxN3jHHz08zhGnqKDSCkkH6SDqKAzRhbwvqw6GI9/c9uuTzfSJg7CTWeNjBhtM9ip2r
XUq3+QDxpQU9KJylWE7ByKjDCe7N15tOK9W6EW3GwlheLqJwaZvwx0qWtAMGd2BfcdXSpWelpFjt
ES6W4cUbHFONEFPgEE43SH00USUQsQvMbnVesVMmHubaLW65pIAy/jj2L4KABAVIZ3VkrqLtLcDD
smseUvnK7OAr3LQ1u86jd4yuAfbn6tG9cWIlpoofGpYEJSVvXZiTyQPFtKmBUptGm7HLDQErFkDN
rAIipob9fgNBSsNgO+5V2PGlPa+Wgs++QWgBCgrDJNUOMr3KJI/mBz435khxDXf4Z8auspQ0UArY
SMkyKyNoghA1EI6kx7AngcziL0g5eJP3nxt4HT7DQItAuMXUpr1acfQC32y4Tl5nGBgyUBSC5XSl
EgJFkcc0xhML70/UUcvfWxyiH30Ohg98/EEKQkK4g8pSSpxINXdshpW1wUbVHf+/V7tUsW+J0CQP
j2oX+WVuF38IsC/K13teYlxKcP7roLkUpH9Ul9Lbn/d7FZuI5vO6SJTs8ZTxGtxgXnprIDrGtQa5
CBMRsezgtMIH66spWVgVZNh8dEP+mxKxkU9zSkEQ6HUTwVCgFYlMnddlvowcZyRD9OYVbUD8eVM4
8YejFCcUzTbWcvYjIEtzZV0MeEP06hsMnvGiXFD736MzE2+IF2z0LsCKjaGlK1smUvhASacuIVTC
gNPuXABiPRTPpigmt3mn40lyc6KxlcmfgBHepWtZJZ1Y3Lm1zVIO9hzuuoGpqpycdbDqf/jdP3jp
jn8JsnR5XcAL6rIPUyUcmTm3CJWr48gd+8r2Uko4mYGYrhJ1x75n6EdtPYPj+B52khrnYVaEDWqV
E9LfsPiuCxaIDpaEE0lRs1NX3Q3V6/n5HdPD9O14g4GltKXZqjFtc9pwzeWja1eDwEwfpW3qG3/5
s6y3bxxsIPRSKw0IFrsb6uqmu+a6JXzYXiK+L2utp8k+H6eMWjKpnnirN4AYln9oRSaERLs30ei9
a6ZAY8O8YPYRp54Go3DMcIaaCAjMwMlrLRPlQ4JsBCgQ5MHNGijQ1+WYNCldbHunCMdQRHrqk8xP
sVaQk3jYP0UghUCMJu1apAUkqddqgch+Ho9FFZFb4O+8CmZXYfxqbRL3OwNsB65dxF93JwN7Vw9S
ry7YzbVIIPEOfS/ktKcnJpvUgOsmowalgCDclM+WAetaPypoGQ8djoVhO1x20gtrGmqNxyOrfNOt
tH76FkAa9kMg3wNY6dwmkIErBxmGXqsbXzYOGIvfe9IaH+SGUNlKZ6eCs+65wQEjVRgwYOsCSKJe
rglY83/O5puYHls3cuyJihCr6uAF0eYus14mWoaVrCAtM+8XN110HQPGPuxAoCSesHVXFdZK9WLa
AD2X26h1qLsrjOrazHl/+ryAYFc36OpADgGZEp0pu3o1Bm5AfoVnpoVWL8/WxdiLnfaNloyHgfMI
CuTVT0sub/EqlokpEy5bXkVGuH61SmqqMVucqp6iaIA1PSA4De06HSdtfw+Zk07uB/Bw6+jNK/2J
8MNld79AnH+Dzo3oEaegox9rKc1xSJMYeZGBp0d0yqshViKVbkfTabiI5swyy/ccfBmA364H4qfo
xr/Tao/M2Ea5aO5C5HNXfBIu16Oak/7HOWjwc44mE0fnIEb/pGSOHRtjQRtgM3hHB2DBqdm4ASaR
WqHlJnHIVx2CtfTsp08++0DvhIVDcfftxFEW5SzjN1Rlz40i/fjLuL4e26VzgnpckvnMZTTpBlys
tF+P79prRrezXnS1TtiPkCtNmO2g1chdwWjL6NnF4eBBQzl0bHn7eWlMVtzoOT7F8CsRmeETxfOK
V1yYf66yqnAQgNsvYRZJQHBwMIDURE0SfBBOyoNzSMRrYAxPclBRptmH/Bn2Y08Qb+MalY4AkOyj
VuJDXfhu/aKvJn2KBm9xT14YMZBS8H6Z9rtWpAVcwX0MX/P4xOq7MS7P/VYhuJE6BOYmKvDOmtee
m558y3sQrO79EtcttB5Wxq+H5g+WLsOirO3u2Bnaid1NVQwS0F/JYQuzceH/Jd/MMubbES2HWrWk
F2KYozfW04CJ8yXhzmjGCYzaE4XcaWW/PKrLuI4aqbbpA/CIoRDYR0X4s0aRJiCvTDumIbll3Di6
am6C6t+RHk0hkdVT1+5hR4ubBZvxPGmhHOCTaf1zBhyG2A5cmddmGrjcb0ushKzYQmpPWrAN8rxy
41odIL8A8DK4kmTeTUqQlA13KO3rplLPaqkqDsQhrR+zdSChT0w9LVILBwjenMV29jacq5J6hkVg
J/JnOEa91IYqU4tH2DGpC43LV2L0CpKmZkEMOCenxG/9ZtwLRLBUYVbcHT8+80VBdWjPKIOoemhD
QmgD+VNch43paCaPscrW2uFlzlkgfAz1hISG6HjRArRv/hHbBSYco1OwHNoafPNQ4ifWErFDxtdX
vR/1euUf77drazbqH+TAmOsseNy+5ef7mP836x3wT4PL/V+fMNEbcDbc3pfdR4DcWsH2J8/t14p7
lM3PDiiUYK9bfpWnHVBWVIx7j0M15Hi6hFwUOEbQD4CBg2NkRPHFO+sK35QaeYiRtwYeRvulujHk
k7NIgF9v2gbEQuhNpVQmN9sSRHkS7WKC5/NGey4hsuk1L0yjRSUXIohjuYwhPRGZuuyag1r/SOpo
dGjaArj6ufBJnr4SRs5BpePtj2B0liUyC6nbcYrF0PFOSvvK/wejRo4elth6uTbvHgGJLqd22lpg
EGhjIJ4+ZksHi0cdb0/oJmhP6xP0n5AWlxltfyFt9tJ7wo5EMGNTietjTPZl5sls0Lkaze6oN6/R
r8DvsQKkugsSUMJPRA/6KQuho55F2igg42S3HS+d1HPGPTtZcPhL9DtzY69e75rYkzwpbcSgxZKV
E56qXWKid4P+cejl0L/PLByOUl6XAIdVeX7jyt/GVS0vda9bTUM+cGuCKM6D368noB1BwFfBXMPZ
3QiUBl/ZqhxKwFqByz+dfTF0YC32bPP3hOyUwy+3UCSzwsZExizwFibIBYTLiZKx5x7OrZLT/5Qi
eO17KiyaNyju2l4wsgVxW+A6ih6ej1GMNkVAhbNVonBulgA2VBJ8Z1MM8hrGJHhkKIGUGrm8SP64
p3GdEJWS79xz9vCM5BLKMXk6950wI/+aIGBXFR+AltjfPJwqnZsOLwjlzUmwmWipZ6ZCFULhyNuT
LyzVQ3fR+P1fsz8Wjj5YTsnON1f7qB13d9KzHQrConsPQIigNHuqREsLOxbG5pu23QkubMaH9YMb
PUEtZMaDFWtA6eX/PAoZ23C6Mx0iRHTm5Ho+WFvc0cR8GDvqNTVC+hHYXcm0QTFBvv2HZ83W/N9j
yJsQDTzGckppFPn4tUYkSxWr4wlI4CclG/a8OiKzCYxlNYaH/DFo9f4/WDPfbo0peuNXbBcULc9D
P23YzeMbuUZKSKDkjp2x0LdefND9WzZULoZJ6odUJINhc06AS9eUx2CFJ0S5XO6ey6jSLO7y7TDM
wQbJs2GDWfMYfPaWfQNJb5TCZP/ooAqD57czZ9fZwmdwqiqjyqOeAU/BLFOZKoSeJfX7gKydknuh
XMgRVWSG/85zRFtcFSxYivWz5A5zxnVI3zY26hxNKIm63x2rS2l0NRCy4kL3SgRAnSCMlUAW4n6y
05ZQkZ1v9EdH8oXI1rmO2cfsWg7mG56xsLdPbdm+xB0dZLXDDsg4euFs8kLj231nWKcJTU3LZo2Z
DUQVLCS5CE9wwcHy+MUa6ir5kbKx3skF/SuoomkcKM/bVuqarGejVLDkWCy3/Qe26UHkQDjoOYB5
cKEF8pc1KpYKD61U0w1HBllz7TPyZmlbEbKDk2BaDt91AH+GpuXXkYPU3Veb3kYGh5ikegaayF96
QVSLfUEMx2OpNGD0ut+DtgSCFvA3mCP6cbXO0pwjYwgzO5GBDjqPey4fElxv3+zVyv+OHZT0Sj9j
HFE23FF1mmeL9YmAyPwwv6D4PsCd8NyIp5EUdHo7sYoyyRL+ARYmouWcf1ckpROtrbS5tF1qww9v
6Ii6Mjl7kukvQuQ1693kB0FrchwyrgRXrLHkN0hDUQBIb1WF8IfiPBgWUftbaWbQpArJ2nnXxchP
YVzzWR+36JH3dc7seMmoQdoGCOEsk99CxtNXLTOHAceH+U+bS9g4sAGWp/mSMdHLqL1nz7rLQAUV
pGUjZ6Pg29CAI3IM3Qwb/JzgxEcw0mym1vfmDNvcyppbBNYZsSoZZPsaFNRiSPkdsxPsdrK3zOUA
2B6wUA+3ahpT6tlkGXeyDTeBc1Sy4D01UJaokL5k+DYT6Px02J2ljJok60IeS1CwFA4BvRDHYu0/
Cm09tjYx/nuaVucZw/nRXtV/CVlw9RIVcU0Mtq3EHvyqt9qRNvg1R0WekaSkjJTT+7mLwR5VXVXw
jdNObCdIrx9Efg5vqydq2CJyNDkW99MhM5MnmDzRsvhWxBxKfBLQ2mFgaa7byWVkdZLVL5kktok2
o4RtWMVShluPBdlbQUoJleYGpLCNKEil/P0oo7f7ojR6N3XqabNKkf54u663oBcS90nTyVirYDYu
u/EY+JQsxD2ztp6LSWmhFHfPcch/xdIty/IXhkbW4syue3B5BL9soBrREcyZhMa733DZJN1XGqbw
XJYT4vEyRJpUL7H4mhoAf4EJhWk+gc8J4b3i5aQx0DyUm37ad2mXbqPrKyR6aRgWbvrxQvx7iMIo
uZ6AkCytmbzGaVrH94/dU1qk/VIpeIsH7W0ArcKRyjL82CdhLPwS7jE9usH5lHIckyDcpr2ZOzuo
AzheOSZag7pxiJDNEI2fXDIpCodvEkA3uosxTns0WyBZa5L2o/wYpqRE0bAkyPHcVPGYirPTSTjt
cQ8GbymTVV9AFpdIWd2aRW8JcI0z2InnEY6aPKU4ODJjvTVXQi/tBnB6me4rDIHHpKfsxh3FNLi0
jIiYqJjmuXQeh5q3FmTqC6hM2cFoXiVUyeBOD468LFgghvxQnYJTW1kwXYThK+biyOR/PDDtuq5W
Sc4ZL5ix5NQXNKgmwvTGbcOYG4bkxVXRYWYSZ/gxLd9bY0V3LXBpsvNesNzIzRbvjk1k8V+oZOUk
PXUF4F3nLwYHGfznaMNE0DvLDhIP9r60CKU8ZTGtqIQ5s1RPJ2vj3Ut4oT3eVdXb7laMZSJj1Sto
MZUV/RiqwPh+MJgH0c8UUEd4nOyxP0xrMZBDifw/ngmgX+ONM971ADeedqOXamDtiHWT+HInQ7fm
h3ndQZQ8FAe+UyLpBlvyKHUGVhqyXsG78lVyDhD9wfmyVFyoczVi7EUjsq015S/Ug4XAtLBiQHhn
MlTRo+FNFDIqkajKbWk72lnJWjv8ZnLdfUX5E1dyEIkA7Uh0JOdYoFrL0qKSFWCmoiB9vw4uHsvZ
sogZMii9XeUknuPd6vJpksJzIXEBZ20zn+qnm8YtFc0UZpHy0PxfE1XY1cjHinR00Fot+hB2QiJT
PrF6+W1OxsLfyxYlJkoJMyoXbjGQ6etf25s8Nzf+tJYO9lsrZhV7fJMv+xbh9/gpcqi5bh8LtYw8
1KP588Jh365Eck8Zd+rPlSr/TSfLcDTRqqjQ1tbeLI6HBtCuwyeJusC1bZPVcEtE6HthMjmw2rqm
yU48xokFgdNJfbB2BQKwweEGClrjFF6nXqehy8A9LsGUZajPaGyqy5kconWwntl4AGCEEyYWPpag
BsSoKAG6B3fqSUljGQ4rnIgzz8e9Rlpszns5lDqaF8CY5V9ARrnN7tDO9qWHj970ZNt1d6U44115
Xil0I4ODsAvaSMDY79tNN0WjRupkbwVoxJxhY5Zo64ATTfEcvVReMM8nmIzxUZ3icd6ioxUwbqdV
y5LeWSAbmNJgvXHeG2SS1wisF9L2IJ+IyHvklZmvjQGYpNM1b5Ycad092DUCxFQhy/YaNTeYnXxJ
wHGgvuMSUtBw8pEjOUH4Jj0yNIIWKzi8YxxITETH2VgM2nsu4QI2Zzet9vdXFkAxCF1S8FQWq10J
vAZN5o1OfOxACXsP6baSgKPR3zRhMScysaQrwWHEeR4kkbvJC7tmAMgKsPf6+JrHdTlVSpLeGj6W
zmNz2oCX0+/2nL4IBMdlOVrprZGFb4XWt5QUaD4D3YO0Yy5xw18I4vISgbHObDc0kBrE3n/VVmjx
OWZ8cNkKAJUlbcV9V8LNkYxi3VCJj2zBi40sUN0yEnG7rIyK6zEaEbQJ5+ZSXCzuMyLAMRfJEV+j
6ZjSGHxwZMW6VoIRLyRorfFWc1LkrUAdIhi0cTVEAzd5eMFbqafbDySZqVSew3mF8IdAmF9gKmyS
hoPxtZSBWi3z7sv/PIVonFfrCgi9sDXEWwbH4h6qmg+Cv6oIC3wTUSvwnAfd6xF3rCzSI/K1OIA/
x1aVTJB+ImKlJzv70nxKMIxWnpgeEfZm3mW9OclLUBItKKu+UVa+U8wvQk7gpX9tnONo12sqf0bL
+SoCu5kDojoCaMxbTOUxAGUYge1ZUH6ILnhkjvsYK/cTL5+/GQg+3oztF5N4+siZLNdC0XtIdAWI
vztstEYsMigcf4Hw81xTGTthw+h+q6b0O80tYxyQG/o7c6tuPTriVQrGAFvMnhL54uvvsrhLv0bn
WoZrA51tcMLYK0dEpSIEo4Jg2JW5QIH6GybswJUfkjwb69268gC7C7yViRWVU3Z/WJFXpVJK32mq
fwhoSTlGZXwJWihv2jtgLivFScNVAj5lIYG5idWC/bJBUrJpLxQQGB78pUDx1DXyvPJPdSdoAqwy
oNrGynth1DPkvEFgj3dlbpdy4Yl5wAdBoOX8l3k46rP6qABoAQHBqs2wPcHJDmswmz3DdgvEDlJp
Lu13O5gLKJLbbuM5QQS2DkJupKSV/y339mI5yL6ib6JpIMcslyvKjDLNinVS8BgSk6+Vk1l6rwrS
UqRzSnLzbVEmVLXjj7JETgLpYwhU2n+GeizzkBiR3Ie67nOLF+hFEpEwdswsGHrDdHCvNKcWW9As
qlarwxxU+XkXzSDHTy6ESpyODfYq7DatCfoMiOddywdSkNHGGdmdq8rHfbNA1AOWpXcoyRD7hC30
CVWHcGgnayNGSehwrkUJR35BI0uXMNzHmqdDbDZTXtpOtuz/29XgeZODNezFnubPDWawG9n+hWTc
7gvgfABm9kUTCyBxp8IW7QOBjvrIb11pP+jrqTaqpfR7cISMgqv0VYc+OKFqiIQX85Ij+FVWbr8s
G5xeIaYRs+diFhUuh68kRqkXUrNVCvqhMNOG1TW2kQf1MtijkAK6+UVlcnKRIWcywUAoxxms+81B
qO9fSrkVP38SppQW+Ss3MFnGhchrUwci5kxAal2YcN0bVVBJZcLSyTKr2dnaVeIeQ8qvKnPFf10f
VqcNPNHADE5qzl22KvXyYckhWaWwbFFd/ZQ9qJFpV3kVyH5xc6aYmnPynD3BoWgYhaRPryJ6SMHc
A8wDjj+cb0taupveODeCTybxip6LfI0qBV2yFUXh1OTQodY0LNjVSBK+AkBVCYdimyzncD8nm/nF
XRez3pP9poGLem4BF7OWZCxXmwssWWefoaXu+yWIc6TSviMXAYXvOQShBWEXJrQjuRrpAmQInkEN
Bu8wUWDMcL2fba3zak8CKK1SeaVVjUGwE5Q2ES+UAJxNqG1vIld/HFoza0inPHj3LjbyrXQMk9Hw
40zKL7Xh91v81n2ACw6/964EXHggk+NyasyylAIo1O8GaAfY2jUHLt+qns8oxHnFKGmCijTPbVx0
/4+j4baER9kbgHQcIGQxIoPli5pmChT8QO0pdlCVCtz9bUMY6GIJ84tp71AlQhhHNmYLnWj/U0tD
IB4BY5oLc9y94Sn9Jycd0OrUXmCr4PM8XlyRbl0lYBUaA76B+cymosu8DZ8yjT/TTWxjT8PAXKwR
hQHCpW1ONJGSzUFO9aw8e8jwU/WjX30zcdvF7F2TgdKSjNZrq5ejamckzcz5wdnSSG0USJafT/a7
DFK3Ta639EG1GpoQzs9NfFbPZGCaIaXE7rsGk9jB7gaJQsFkydS6hbS1F7TXTWMyB9CbaN6+6BBY
jOM+imdlMILtVfkxc2nd9ebttPPvPo/tBVPTSOhVXzhUPb3xY6w4rQ5GMWk+hdt2QfYKLYEmwqwB
Ryobdcy4e/00UOv2AHzvKASp3LfEByU0W304CI1Qfz5jpdP42jAOZWX2Ay0YXgK53xtWAyaVtXfr
X9th5aqZwR0Fxw9Vcv2FmA4Gh3Hv73eC13Ni/bdjg+9ttsIfZLkCkKqW16rbrZKWuVSitoKnubbS
l5jbTMO3Sm1UNHabL1g13+9zcVukDRTELrDvfbdQ55wuM/7Y2sQBPbzt+oAK1wNvVaFBeShk0/Dh
gXzpIfeSQi0yXQRSRAyaBpnuFUMryyKPo91qKDSGtwUkeJFbmMIvh8yHZqjgd68M+96/KJuRsZnw
na3xC7rDFCmysfMRxZodJ5MNpGx829aivtFtybcqPH0RcpIGw4XOhPWSHUb3wHbbPffhrUZA1+zz
oGH4laYnBZK+ip0BzMDx+XjoB53X51+ATeOZZNlM2zGzrCXpC/ox7bKPjTrfB1Pz0ydurm3gx61e
3JrfY1GnObWXPbkum/IFy+Lv5oQc/X1FsOZKvEPKAmg3OmlfAS+3kUBSkx8qMrdKgAodvSrFA9kf
fs5tnmx3ogg4UUpjXIKga7RPWkAwwsh5R/q7P/AUdcTjW/LZ8j9BzpzrJYGYbgx5QK0cG3VXbsOD
zhv2yQmt1QLHtvkZpGioUdhyVhgbi/2CRV0vKLY79dVlAbRK93VNyHDn3VJ8KaKBk7Th/g52PBPc
E0JVH1aAi2Ol8uWyAfksmwYJQR7t0knDHhclKhvFIuHVRAZmTgiWoH/zBtv6ETNPIQiKPw3I9A54
A/11Yw7i/EUr5OW5vQW9ObJy/3Ab+AC2vZSdnkkUjbsUwaV/+hur5kQChZs58l3roN0bhl3pLMZP
G0tfLfaXFpJISer5YurhoMMw+Bi2wR8j4fiEjkJYJP0CGmma1gL4mr9nc0XDuSySUJUNp+1Ah+xl
cTejETRJm/9DTBZVGv/FZiAk9Mo0+F8kHJ211k+mJFvFFxXGjCgrYVvlhI71zk8MVer/rqu1Xovd
4ntiTjTDaQMt9k1OAzsoa4qgtLmPJjEEszToh6IcWrthOoZdBn2+VxLLy850ZZft+rS51GUAVAo9
oqeIK2JkWdUHqzyxp99unhsrx/z966rA0uQP3Htjiw2DemTOp0DZyCdWFPb7hNEBSTUJweFHgpnG
dy7Y+5MAWEWEqbPLa7/eUNbIyACVgMFuzbJnPE9/SSfIUBQPndrKzTGRi2FIuQgy4j5dZ0vaRh1U
v/OTQg/FIBT60zrI1sG/f8DVdwbNdxFUJsattbRAPnxjGJjuincampD8uR3eCHrKUOs1PTuKx9JQ
zJDHKStil9AOOLqtwNc0cy9gUjRtVRe0+exNX9BLVBn1KDabhOoRPPEQsmyGczpBTIjviYJ1ku8o
BVNJtBXHSVbzZ5wGIr5pi+GtPRLFLdzacg9FZeoC79qoBTxqcftrVSYuMC0yowaep15ZuecfpCAA
pad2tw7101so5TX3H4DZkEfRiSVG+xaqwB7/hezZ0vUBPkXQfIeEWeiDDO2ffydqsL5GvWb/o221
4wCKalFWm2GxyMJ+ohCOfleGEluVWO8uvLPd29/dEivGEFJGlS6EGppVLQyMnlUvFw+3Q07/L6nO
9zPkLoFJURTJejduVVVLEJu+9SYD3vq5wwsSav7q7lWUKXbSIY4xhNKrhyDb/8fWNzxyIygLi1sD
WfwOBU56tu0wV5IT5tHeWlsGn+ilvtZ4JNypjn+VuPGzIcx5ShlXk/pPJpPh04xQdT3EHAEkuW0Q
YN7j6hUR2Zn7Z2Jyvt0rDCUXJ2BEJXhfIwoPpKkq0IfXBSaPN7OO//Qep64WiVIuVYLX+BItLxjh
PONycJScNetwqlzBITTRCUuqKnvWqChXfUQ3TQh0C3bsNbaVTo5RMLOdleUsRMnzXYTJiIoZcb4m
u8BGMWSdWRtpoT+xeBpKN1uup4g4KGaVKde37cuF8uJUK9/uZmDYUaBV9m/eocF4B2htK7se3lRA
/m7RpUUtXs7kytsKy3pMVGfqQZXHEtL+Gr8gD3+IPH52RsJJhC07tiHun33WBYfkZ50RTOGEb6V/
Pfln8jUPDJOA6S0tdAqspbtmRhD+P2JcsKl5sgW8Yxwv7JelUsUJZVTwOk/HQ5orM46dsvaVfDgo
vre+qJhTU/0IKFNlIutQ2k2DutMujH5Loci145oQFjqwh+oOnekF7p+CtQZQhdZbRX+VTDgL97jC
EtbYMp937aF0QCnhU8to+cBbjfvfIrKE6VM9+Tw+sZbqx5T5OwvheX51NBbasx9fVSkG1aPlxsop
5JTpDGN8x5C6audyojDzK+WxHBbfUeEdnSNBikU9wbC73byDKgaYXa1vnox2HP8o7KAKqPLn/Ey2
+SFBLZBI8EGI9XNtfcPcZi6avPIoTCjqz8MMplt2FSCYAK8mfRashltm4OHQS6nn4hYysSwcflA6
7kwFWe8+bd/mCPDkbkgK+zugj6nIoqQzUwglG+EANXFDu0UjcauuzOG1iP9oZYhEENKKa12EY6hl
11zFopMK89qJMVyyAtLoS6mVY07fQ5/vLpSVPa37r8ChQ6XkN0jk7Z7WtJfygYuftZR/b5flJEad
haztaz06aoAvvtBPN8lLZtzw37+/e6oeiJeNbZhW7oYjMNVzZn/a3+VWqHUQjQ4FGtuuNDt2fvMi
WOim81+xpXl0K3n8fX0w5QQVnG+JWLQaECe3ri9FCsSjGg4rb5mJqR+/hj1HqUXzgJvbuSvXzDn+
GwTSjO1iALt3aXqnJBf/MZHDEKRp8GOy1rXpxvLoS8olKVZg+7BHCHTFdb5C0Ky6O3uQNL1bYQ76
xfMD0xM6ntrPpClAI4wACx2U7sde1S75jCGhbNnF5BSEXpLHYRaHc5IL/3tiHT184MUxihI4/kou
H9LbkRU1THgAJF8rbC5HYACZfHhZA44CuyybLt/3O5ScTBe4bCH4Mjy/yh7Pn22LzHkBqqp5hp9G
JOA5CkErHI86LrcWXF3WnXHp5JSLKttQNjZPjv4o0o9qSypBL1qa2dO9KnAuv8+rB3ExN8mSaF3q
fhBlAWanbM3gC8roomlVTVUW5BtzShzhLlknKRkie7T6BHstBmftldu66dhdQPQrSnS2Ugyk348r
878yY57gS7JB8oJHaUPEgepiS/bNW5qS2rA7gf2rKJ9IloCEKJclnQV/u5TvSFcei5/5gI3hB/LY
cDXB4I11dXiVQD3MT406bzCrTcz5DC5YB2U0oJ+YukqcLfDZsctnqr45kESM2XPvWeKq/2Hlua0q
TyNopZ6CGLlV5ojH/4yz3vhGIqIeKzYBBd0Z8WCAlhBbDjGKRBDO9J8p7r3psgrMLqW8dLDhRBlv
4wM/x0CUADIZhcCjn9S2um2Jaotu9JNvYkYXd1cd/fcJiiyvRQz8UEqZzVUWV7adxjY1YggpdhsP
x/dW3X+vXZeeoaZ2P5wlhrkqpWdrnQKA3KOJxlHEwct+kuoOKkCwz078TxeD1Z2roFzEs3IoqXF7
004oCfxDL7V3AUzcUy2neKf3ClJ6abGP8XjQM6m1sULgWJmTcdj1R8yYVkb8LiZXP+yFd94cw0rI
79DlB7Ogt+nXEftEsFIAPTLRqc+bmjjXOBbV8LNufdMqs+2daXz2lFt55NtBquZwNOGuAoEPgNqj
uc4kk2GKuEGTr7yoP4hphgNQ0EDZUMTsk6E/lNkPHArl3SIbiZMBstMNoTv8nRQe7rziU6O7nUi6
8voSln6tKbYAXUCdmKF/cZoknQFbMwsl1/BImvpPVfvSCJfd6SXVAkZOnBanVhTmgLH9r28hR8yF
2F8yDuRGJbRYbM/4tbMkh12XmQa8WzIz4mSvhWuaWK7Qv/lzdfpeqV4a3Qk7DbNd1uqAh5Efi9mo
EwWy57t1M7SbNH7q/39Rmlk9A0FE4/SfkkU9hXIfNI9r1JpAQRcTi/+wGqbGmwCDCGae5zVdyOIi
OMbfMCOpicmCbV/Y6wX31Q9KfoTui+KOSUMzENM6HcFJeVKMvD2V87krfxCxeqIdtXJxZc3/tGkp
EHXynyCtDzi/2UOdfRsm2qSD++Gtkr0VbBnaMchOHH9J6OGeIH6/4sq5FJpXDba2PlhI24rt0A4O
aEA7YeTKGB8MpXWCPMNUWqoWq7O+Mf4fTKoJbTxU0VboZnr9O3ChRphOSIK+LBver/LJft4Hrwm4
Paw0ZtCY+CrMaBFEURfSldQr2ONZOg7Ww6eqpJP1Ff1Al32whca9VwnaN6VAltyNNaeAD2H37OpM
Ai43maEkAahxjiFOuVbHLhqJM4laDthPZ94tAIf+TOUnN4Myklx3rXjuK3Ksw3iWpy0RiSLaFN94
iaIBQ9EoEgOwPGJAWjCSZ9hbk5TwzpGt/kLUYqZNM1kQL/U91K40MUqosYZIzNvqb8WixEJUAWSf
yV/0sO/3wcJlWblWUz8g/OgQ/zJTYk5GQNkrQtIdzl4GcxTHY1gcBGG4g0iSrYlRIQ5EVdGm3YoJ
vpvZEApURYMGmd2yzKrL7qtjnviEntvr2j7QcLVMyg9doBMlZcQR09XhcX4qnVz1YY+LAPqVDM+6
WNz3OUtrhf+nnCJsgVtdvHZZu6ondfhzPfZ3XqCUiq/hsBVAJQsYhT4jHU/PR3qmoK3VT+QJirOi
m9FicUir7Dt3AhvWud34S/HyiEdrvnsj2aI3m0nJMlrPFaebjGf4GEzGqEAMLkawB4ILewXRZKAN
isz+en0V2sqAazRPebd6S/1pqdBOuPJpY3Wec16BFhACnvFuneN4pt3HPl2n71Y0mlSwcipPutoG
5qs4XsUDSx0hfAfKkGU4nIAojYmdEdwYocp1f6aLvwAkcvq8QMjJKPXGB70WyGqyb36tRwNv7u2q
byf5RNcEAqrq7VEfvWZ8PwcqRk82LTB+JZkZYGfGpZJ+sJDfBgdIBy5PvvqcRfdXzdEss/HJyLVe
reWnEBZjD0mrFZLnpmxkJ6N6KQHIv/J+Ou9b14SyU3I5E7Xy2k0cYcMhyzWY8n1ZlOacRB1R/QS0
JhbKHL57E/JGmoGAAmPp6I4bw82GOvD2w/NIDdeyboxX0/+9s/03OE9TT27HqBDSYe8gYlJu6B7M
a1H2wYbvA/iYoqtuB+aKk+GtOoaeGyaf2fBTNrx1c89aXTXvwuUjyfmPRxTlv6Kab/FkEkQ09HEA
k8qptFIrTAEbklX/GPAgNC/0Bgm5unFcqJfJUX1ayUkdwwexTsyvTWI3Xbh0xpETMGy+oGbjrpHz
P5VGXxfKVteypOuT5ky5jgKOp88z2k5vk+LwmBCN7z/uiu5EJY0JTTumNmM+OZ+miBquAR1XFdiF
0c5vuD4ZGJ3saHARsYXOwqhY/Q918Z/fU2XgMa6XRg/nA+eRyT2f84G52N+noF07PaKVm2Sn9i/0
dVgjFhiNpb7mmo/7ZoaLniuvv14KNOru8w8EpEXnxqpFsYGg0Ai2xMP2hL29Xd40QSL3T3ceTZon
oxGt6AShO79dClp9SEYStvX5AeA02/5FtQtk/O/S9MAO90D2gzGadI4NVNxfbcRHyfy1ELCLZ54E
CokC6831M7UZv8Wtfkw/S1hzaloYVBIh7+XslmxPi6FI/cer+p/C7VoEUDFzIhUtiaYx5Y+uPuX4
XnClYkg9IA7gyiJaDp0WEIIUFvXo1NiIJYNenCsBmRcG5IAT08wSR9QH089+d5gnzQw67JL46/su
sm/FRFbvbv3+m6FCC6rcDrS9CSGdDQIZLPK/olipd5XN+Cj0xNDRrbFu2bnijgpJqNFqGI08M0eb
cjLczfIV0odLWES0ni0aKJVuulwYfzYHcqp+mnU0qN9/15u7xVlSM1xT4nAkxajSYSHr4fWtKEVV
vIS/ho5VZwmnIFA5JHi2ifC/DKR/cd8GS7uu7rAS8+jeCwQsOOTojQFO2sFSz0ZC6PA3CJrPH4/D
uIG1vhwt/oqgWLsjotb3ku1MYp5u/kgN6IDDdqtvwZa5A6FI4tlXcYVjkSsDlELQ19ochmHiFkcc
3kitRslmx7rZe/Ve311V4hZhLLl6Nxxlx+KRZ8Rdz3DaoYE83GG75cu8KQENBFxd0GUE8wAzC4pQ
MKi9p5vP8IaZUmzEWj87YTADp4BCUI8HUnkgR9RMzCvBN0FbTeWZk6bOstg6v1Ih4kfNKR3TiiBa
nUhG+Fqhod/CwXrVOQoWXrqNZrCkc2BaJPPluSaHZcm/OyFbnsDF4/4fDtEDxtyWTta/ymiSKxSE
xofIL9GNmHi4dvlkxKqqiO/aJ4wsbAT+AThmH1RUKhTD+tssa5JyunUVRAijwMi7OpczxpaImRse
CjgHyudc1xrvAO/F4CamPO7DbYZu22MWaNTxO4wCAxRjrUHEAtVvmLKNOKxX162jYLarJoyvMzz6
DT/kcNMpTQS+qiHexfnJmsXgGU5RYEsbQbtJ0cDPq/A4rpEoSgAazVSXx1itSm+9wTpivCYpE5i3
zejUzibpOtFPUDP/QFOHe8VSD+z4pRL4EsOJ2x5BE2wYXGzq8S4QoAD6PHNmDiK3KWbndp+E/1+F
NZd5OB15nNuiFVWaFBzj1zQomfvVKXxBPTYK6in96vUQlc5+htkW+gPO0KA5JlKwgHlyDh1pPP24
uoee3HHNyC4zZRVA7AuQyaGqpM9VDVxoMICOwC6vL0UAZR7XdW3MiQokvEF26Kah0VXeTHQzFGCc
1Fx4hi+bTgtzOZ22LB3R0zlyR12yrEXmZFDPm8EOwTMwjcmUtgatEaIeRsuyBZ/TRnTGfqnQJLN6
7AuYoo8sDsmjtPF9xwyjBTk9WAj1w2m0XsdW8wp9EM8AzGCZhi14nLdHmRZt9qyuTeHzSnUJ8kJ1
k1xYy2um6IiZJPsZMxTg9fpTsmyVIoU4S6JB0cYUOo63Nvvs5iNDO035KZCBqxxVqr+sGEB2p5ex
tJctvHc7oV5xnW6/FXYSD6C2sFzSkV4KkGa7oKuHHcJgaYxYMz1xnKClOR9pMBZprsHaR2gVeTPY
+O8LughPlFRXpjiJB7LY17SNEUQ82sLPh3yMqlQfffS89eT2t1spdtVEOOdfmmzp1j8fiogPRPuF
Hs+vKbGMTqqapqYQBylPdj1byHf8tI93NKCOrNOt20imaMhaxRLHDlOkdcXUWgiZSb//xQQx0td7
bH7aCL2Bc4tP0pmUU7cxHjVn7N68Dya3GlN3ltLW2XTRbOvlodaEV9UPRpyW4yEx5UqXgq2tfyq+
aB9UlbPc/LAgYVDgG/bjQaw0VaShG9/rY+pzI7zNwTO/x27lxdDeAtR/o8yRC2AOlTW2iRzGPoeH
AKF9ZTJz8qFfBpaKLZLWLSHZbDaf9hMExeLeZzRg39LYjUaAWlDLfaSQYigJ3j6KVomDE1dXe93l
d0QJpjgOZRAEyJSPh3dRTYe0pe7WH3u35GmpbZeYKAmsbDeDKOTKIyGHLye2BCRzE6jvjm3AmL/C
wFMGzPj7hHCaUdc14MXbheplqrnDpf/yPigE+HvqY/ag8Ij4skBHuwqGyyf/WpsJbGvB5OYgfd3R
d9oBBDV9rMQ/r3FCqIzjID3q/ZR6h3ePVMGJdozphY363Ih3v/aCwncb4U/8nb8cgtIg0E/e1ZHM
90P+J5smJzhAmeURNHYYNKlBf+wrsRo++V8gRDUBw7+1ClB5m4mQ2gywWQCj9UfrA6JiI6GGMHOa
WMqtH2rKiaizo+EVrE25w+zQDaAellTXYo8URr2Cy2tVhMtJBQWSkmBUxCGsSNja0Guay7/4+Rsu
wR4kmoEeSM3ksX//kFJ/AKhdUopzHzVkZJS389sa/VlILELvGb0E2VSs5PM96yHeY3kTyh/V89GS
TT+Fmcy5f3iWG7uWbuYIDlrI9bzNz1lJPhCO2QVhASM64Qe8WqrqixLVrJwRyd+QJdqgRYwg68Wb
gZly64WhhN2e354Z4fBziTzSpt4pv+CYJJlbfJB20og/lTWcL1YpDHqUXEHDE9vjzyETVyDGkWm5
ccL5a2GoyJ7m24Pj9QFVeYI0lxWkpV/45p6o7PNLInLbYezCD02ZIkBx8B+926YtMTCI8HIFr8V1
evZn9elA6l28aE8L9HD2fs1OADSNTSKgd1AfMgwj4E2jlZN+B0b/F8Xw8MDXiz/utTXqWiQGvVpD
0CT6b96DEs135DTVehy+zT8OXEbZDKewdMqLv5bQWVIkbXiTV1Yw830OwomM9y1vkr0Iahl+KcSc
WBBVS/xfqOkekCBrDpqYx3+vw0Wi1F7azXOo3HYsj63FsnWMmpn30VMIycXLA7BdIwQu3KG9yjnP
iOgDKA9PCbsHoUxgpdZx75mv1z3/Qc6HnsWKMKjP+VikNTTkE0zEu0TcBDl6bY+ciFn+SDOi3gWX
h0p6Su+2q95ud6Yppweka4nZH2g6sDeSpj5/mf0hYkPaMwdT3rjukjIWlTTmVw8d6UJ9qExLLcrI
0dKyX89gVAptvz2fWMuBhJtwXJiKifbGNvKyOkMJUknquq0Mk2J0BIy5wukok/jkfNgt5O0rJNvv
l2SrAr3ujiiOpYNEl27CzUNnFNNHZF92xrRFTgV6YpnuXPlSqPdO1HAuqfQLD6M6Ov7P1F9tVlBY
Pp75ETmTYJMmjZyFyxcALUkXz7AheUhI0f2f626T5LoH4AMw8ZFAP2KATIak6vraQQiC+oXYzYoi
4KInHv4+frOOeChX95zwsbwZf1tUa6rzP2hbP+9VYYkcC9GTnEaWnRH4cMRP+cWw2b+e46fXa6K6
jave14WN98BwfqtV5Z2LP8O6Z+PUZVMDLaXs8oXe3RO/BCrs/9EWi3V8SODQWfZufNRpz/6D16C/
EYigWBAg2/kH+RDvQD+EfJcCVAA6UiqUr+hK+XV+YfPC1QUguAr3KBJ/+/7gX74xotxLXTxwLie0
4VqseiY+tO/qiIjwHz0wbeq1iEbatP0cgvDm9DrPQ1wdNXtZTdae4//OHCH15PaC6wBhXkjnW1pl
JHHAlSzwbecTh/9n7ZFcddQqKtkthrU1o3AgcKOKOmsGGVGgSXTlTxUr1Voml10ekedZY3OaH4If
w2B3r1ERWGzk/G/s+8iIznIlYbhJZu4PSTbDyFjx49iudfN8ohndgf4sQovCjjmpiCI+snIkt/0o
TDnOUoCtVCfQUm33FUBvGOou0Eqbf6qLdV1oHAM2XMgT1S5Wfd4xjco9tVYMbawaPZ0cAtjz3Ild
+hjQor8d76JRwiTXH8ADXDjv5opPSSeI6i4qsl1E/ekBgzUs4IKrleBL0030+W+DdinfYX/OFWUK
8ly5jeSAF1IJ8uqwkdc3XwX1nlALiWnp6/fBas0nCXurMiL8ktNhikQOd95P3WNkJSL03k0NYRuo
Xuf/LYezJIrKhtV4nCUuMaUbq095W7zQbUQiN5BUlTkwoHFv8+iAzI0sMNe5Jbo+zSktP6/UIxz4
2hpg/rUM2di6o2dLkC2w9bRiTBd8j96Gn20lglMc2LJkQlIUPMEa6lC/tS8u45YwYrhI0fTQITsT
xTivVKjgK6XDZK/Su1Jloxv9RmCboO5Qu4PU/NDXjW8Q3Tv6/18RESwFMkJzEO91QKL/2E/H2f/2
I1I6/6xhI/QR9+FWZ1/OKzNMqxaRGS1RT5Pxn0vvL/hI4dljY/m6Ji3EgorIc+HWBcuInQcLSA3T
FvoVmCLtxoe2jGZNlbybEiSTImHfShmRigbxlAb1skwlnz2QcFbEE7HWyyAJxmF9fT+o/z+7333h
LYaFxi2k/wjHB5aKnUE51JLzEqCxrjPij5nPuvkVldfnl+HMHoKa9gGzRlcGt+L+8QWFkT4EqC14
apVD/0yKVpBAUbSyNueKcWLaB/YvkJGv8pNVenKvQTXjgmwPXQQPWX1fJZT7aZfUjLFesPqYEOEO
5ahv8OA/t+xBdjdY6RG4t4Vn4bR2w5xHYXEaJTh0dkxjG+3ZiZFUngBwV+CqZayg9/BIHbh0iZMT
8vOyDmTt130pylFnddWPZYpWxZ9d1X3Ch+urNJ+f1sNB+nupOnFEN8nesm2ju1Y4kWXstH7fx5vd
fmuyVBa5CJ4oRyDA55qC/eJxC2SzSA+PE11XwG8POYIP+HxqvSxw3OfICpYhyHIDFHKdNHfr7V0b
04pLBSw6QK5GRWbDKAZLZOF7SujgRCX3nUAgssOLgKTKbnj9sIPHhqlUxyuo/9BEidFtZhJ41BK5
PkddOk14lGbS2EYCLSJPTLEMy3XsSwGr00k58TmJIgoZ58u/DRtYnAFenfABQenqwl88s/6aCo8C
3jM6J92i++9DOfsweXNi6F94IIU1PIYea/wUN9fWFdz0Pk1QoszRfz+QAZgqEqfpVutB8FezyOAD
jZ17aP2eDjA1MQE9+ca92JEJ0aadSaDL0YsE5rlkRY/4I7VeBKC27xAz9mT3Rmeo9Qt8pwNSxqqz
5gFAF3XS7EKwK5gQdwByIkqqrS4HSWN/xxvlFsjohnmI/bpxmYiB9bofHvGS1VsMO5iFnxJj81ps
2MponoyTyf/2oV22YNN6s0X+cEtbInc/jy561IGHKsvM/iuzwtZ5vBSjAc6e6eSd7nkJoGCMEHTJ
DIqcQ/BJm/USxOi5Iaxf44xfc1UhfdlfDWo/FdT01J1Lm745Np4UuwN33wn+2N9iCCIoxEeiERsx
ItMytTFTW8StueQzn4JzgAOSCe/peiFz5yqd6RqdbX3OMVM+spgsNOYpEAQWqOy7eQp/pU75OTtu
Em4Ebd8GclZnh5BBnENJM5ODMUUqWdH/AWYAR98wfqULeC7VCKxr0MekvaAnAcar5iUMVpoPM+WF
OXLf4Ziqih45KddqLQAIqWycO9g6LB6DaJNmEiJqjkSV5z6Sk1AAEtM8i17wvNAUkJ33TNwt5EHi
lnRX3szveCzGZDPH/V40OGGe08nN3gf5inIb09V0ZREgg0BSb0BPUCIVZm+L6+GG68Dqlw+iwbgd
nc2tf9xuv0p1keai1Czf8rCKa3E37zWwCEwKxZ36OWshbPuP7mpx20wT98T1RWN/5LXrSLmDsK8t
3xOAYD/44Y2qIrKsh0IRZNffhUU3I99cUwHhhjOq60hRLXWAyJpUy5+ikeF0Z3Z+gOmZRoZhf8AR
1TxrZbNzS7vzUnSN/mXDH5C6kDeZJKIXSCkkx20CwN1V7XBp/aEC4xx7NvDGKcAjhWv/yQJ6PgK7
FW2945XgI768HTUOWPVZ1hyPa5qV3a0JncqjnXxoylARr3nmAtF1k3g/Nlb2YgaXvH3qdLeMev5L
yWq9LAVorrwI5VaJEcQMTgTmXyLLsS/Wavj6HX0TIlOMyF8vp1CZtAEXlFCUFATC7Lc6z0dPCu8I
okIOFQy6Es7d+SygBfm3aj0+ZSPba1hlzY+8OA+xIo+2Dp473K+xh6ulLfFRaRKmIPMUweztanCp
rgCfVKgkX4C9kNeTG9HKFFioYW8K+AGrADG+OTUMUrdjkbXFwj7ztQrLSFKc5mVPA6JytrdVrdgh
poQOXmJPDSnojnLt7Eo5HBIiI9BpPAOvLcc5ndq7QotfxsBGU1k8WjZYjYHEO4DOqXl6fvfKvU+U
pjna9CwMlpnzH1Xz1XXyYrxen89Ii2Hjy/DXY5BhpNz50FuGHbnsWfU6clLQD/UG+ZEFbnmt6O3n
PofAcgN7YY5I3FvsY9BP21YpDAcTTXB7rM3T17YUu7Avj4o8y66aRyQFe0AdamQ23ctnq6XU0yuq
G3yaqyMXMUoONsJp5AzGG4QCifTlRQ4C4z4qkRSXOWvNe2fWxlFcwOGjWsnwHB57RZKBzrZgrttN
7WNBpAOw6K+7hciEZQUvzxTe8YjVMm+tk1hm2QfnlA3MajYkRx1RSjdK7lS/B9oXb2u33tprk4Bc
nxboeXO2TUPoKVkWW/1cBHYltyXQi4DDfAsY0wIB4T3iGAsfhg3BhU6EpFQ75rLk5LL5hwg9yWVA
+9cE5kskwQLzF1t7KcwmHJ4VXxlISy77vkODMJqD2qfTtKkFkGegEZDNWvfScnunzlComBO3v4m1
Pa6W8oU3xEtgf+8r0Fkvza6FG9ZQVYPlUsdGN8EF6lS2K+SAZahVKix9gaPL/O2cO/gWcZ4o4K53
tWKdfAy4BSpmY3JDT9p60vSmoa6ph/KIqdMRi3v2arhZY7N9lXrFmxSetqB71yK3+L+N16yqoPAa
+xSO1k3mtxNPMioCS7ObgDyvNuAnO/3fbfh0Sq1sSGU4Balgq7agACK1TvpeldFrf8QlXDrmDhOG
3QfW4+Zz+zI+q1zxKjZBeTgnuzl89vRXXTClvN/y8oUv7fzqASlGCIQFj6dJ4wFWS5UiQsj/pZut
h4JmTSjjBO9cfTo7bVzF3/lfBGj6fTvU6AJ6ML51WXd2lTh2BpzT1x6YM6iAfhZCMxN2JhxhJsSP
Bwv5wM+u14Mo4EWxTPBNFM4LFT1ulZoFaxbcaK3ki3RIxaRmUaAGvDaR4qEp7TkGlhurNOWCswzM
mIRJGMBBXvvQAbThOVXgLS0UOnZsX3FtUtqWMp5MOgNVJWtX67R7PYZ8GPXFm8QR2VLhUCFB28yh
ZXJtLsbxLCbTEwMJoI+qCpylV9ji8osH5fEkh0Mf3Ud1AYYgYYFbeWYG7SfL6037tlNfCobT804I
4yaq204OXoT+0bPSEzQNXf0lAD0lqtLVMLcS1muB8Q5x2EwRulPc4+Oj+REuPGo6lxTiZIitBTsz
3WZePepvN9KKtxo4B3pmhR9k3mfzioOtSL/XgUvn1hPVhCpP1mwfn6nNcOWe23pF666DpCJExVjF
JTWGzDV1FzYl1uf22dcPYm7TxI8q4sD025A0M+dr6H7vG8CzSohIbwIr69quPqiTDst5KI6blSJj
UN03BoLwu9xDKSEM5jFI/pbrNrxz0Os9Zq8lV2wsCAQrqS+amhUKD92Yx9qDkyeTYAyeIZOR+ycl
hWrAHNy7ZyF4hTolwnVgNCXLmw75AOW9teBROkztT2+mqnWLaMemYiiueG8m3Im0t/qmgHct3LLu
vTodEXoi6yJneKeN5GrhjS9+m/dh1KRNnCum6cXjPGkN23MaWKOYezlmKeFj03iyZRq/tFKKFNw+
WaiHUyuPJKsVNM2vrA2Zk68dEnknJshcPFXm3htDLGI/S3kCwhRe2TJMeKSz+quEtie/M/HGUlqm
eh/Xr8I7SJ6ei2HDg3FJv9FihiX8YQhIeH1qvZ6q9Kseb3faH8hzwwgFplad0UmGKwC2cFQPLsaq
xKw9xvgamaDe7OuapO1ZqeDE35UakPo9NWh/5Jc7HtULBjLRMccfp4q7TEm45xSBUWDHR7TEIhwp
3EF8FXdWGi9AG8JcZ49z2Rfa9fJXOD8IoqCFQzFFGxfMgJVc81fAqq05Og06DFVh4yNVJ+udCKMs
xFtep85RKTI+nXbbKWiI2zG3d3+8ofRgfL3g39zBvQCfqjAeZshfcuIdr6nav+CoptowP5dBExl/
CbkInRlB6YLdwUdx+n1+udk7mvCExR4HIY1yfQAf34mLcpN1UJ0zUDy8CWT20SlWyIi0b8J1RfZh
xXBjyGpUyA1+asAs7yJhEDD9oM2f8DPLRWLfQAX94bPOa7KFQg65NMeDKeBbJZ9PFrnPzDviRJpM
s2v/flXvekN0YaYQV867pQ5CIhvCnvaBCnA03nV7VnNYoQsjBN894jJlX7jj5JeRAbDwZZ0DpuSb
UDblQy1tjIjcdU71wg/o6OM6ZzXGdrmA/DEr0eUUsDLRMoVyYXQZjDeXYg6XOkqn6xypDFDooXWs
F6uyZj7C0z73xKchvodo343Nkt/1MAZ/OvxZgMSdqv1IxVBgeHITtQQPGHCNmA82SB8kNWU4gk5D
QHx6ilTpoTQQUV4bqsoxtcHfDXCF0j/pG2ymDw/XTRe7FFVcUUZxQRLO0Q4BKphkJjd3SU+NKx2L
Tl8vt4i1nHBgop59+3pyCwBU6OcxoA5CGtLY3ZO96TLGP+2kSDaPPy7tWkTXghd2lPCWvqgF7JIn
27EXqGH8b26y035eFyf9HziWIaWlI19plXJxS0j8eRcI0//yzYqen+aaWXy6U99kZgevM1uchkxX
NnAdNxrGQ7uemGQ6A/y/qWLk7BV4KQBa+Z25uNyTvI2Q6xGvyZ34ZbxvWt+brTaqQ4kB+u7Vh/uo
KgYnVvIGtu69oNmGwInKXFY3cZH4FnCKMfwGI5FN6ZB6ito0omFhnwYIz6QKPnbZ8bCyP8iikJLM
3spRwRoRjkLCfQLkNOz7jONhYxW61NHB7khfMEcgJ4l84poDTeDZ1x2JHIzfTzUgE9ymt0CujXq5
axRBFLgSIMG1I12ib24hkMNCHbsbRp0HXo13Eyg9Ok8ysP73GzG32xN1FXSO6tUK0TQAhz6slhrd
ksuyvYB0wG1KZAHVvIHlNfioSr/iFW6xlbnTC+CdPR6kZKbp59AETYM6bo4OkTgZmfGwSQyMuUJA
Ya4cSIq+TjaBeGXmewdBTcUxSh/n2/ik/VowECXErz+UpBP7ucFw40yb/qTc3ak9jaZROIWbRWNT
crqTqUpsG3uxR7ENHRRseHBYsU/yvcNj43UPqG55MmO94y/RXkS8h1DoLp48mdsqILBk6HCL6aUO
ZZcj2hqAf8ZWtZBCLqgE/0Pd820/ke9uS2LGVi15thmEEYPj2IUEdeZs4rRFm+xC/bPnETdSNo/g
EWXEVl/WL3NOpRAf4Ro4krkN5ulXsWfzrZyVqQ68kMfAgQCH8iYmReUtZONZULcXA1vhSuF74eXo
l96O5it/D5XC0q417MCpX4ofCK91sGdMCtUNsrqDGF8O0P2G8xzR33NrTgtAhEkXQTYPB02b3Jf+
QQqOyLcL2bmnP9eWcRUgyWLA/xvG3DsB8XatELIMKmf9D/EXc8CSmgZxPH+dm9Bu9QaJJqGc/F0i
lGfqQ7IeAkKnJyqqkR9TRAF7AJjY5UPJIHJTKdlgvbzUBNhDkDGS5Ym4NMQBXtrgddr09dvNKlxb
DDX0CcG1s7++B/X1NnufeuhRlY21V//G7De8InjwwDctagMSG9vlG26j11Cd6NopBo1kXzkoE3ST
xj1ogHXtkqqA37jx5sv3pZFVsl9qkYuH2x5ADMWuS3rMURdBu7DfJ2gIH/QvJv9YKskfaOqwEAkw
4kQsswWpn3IpF++J5KMBATkrcKAF9mo1Qno8mRLthsAzpzPpOB3liFqqwjzQ8auAda1NinTP/cVN
dzowmZ2Uj8fKLEXc4nj1rgr+MddMHV7Uyo/vTXDYjpFxHqP9aAI0R4oD7dAmwNJAhZEeDwj7eJ3c
Kj6FzSW191InQxAJ1/ZHU58s3eS8lo8TwyHuPYdr0bKiAf7DRQbf8BaNOLKWddIkohKlMORKmonm
7/C6mrueo5GoyNNPF4CDkWcshZ1ijbbDCUXPv0NXlJ24WTt1sns6ITr/xtdBgiixnjtWGn4loXcq
lzMZ5L0feGjqlhoosgqu5gOg4/rZ07t0UOgnayeDSOnEuBL09zEGm8zNPNmf5jB1My3eE5bQVD4r
WY13IOzfove+uM/ApiSIkED/wF+x4dObJ4s2Pd/j/bVDkdSNY/lzJ/DuzmtkIQKfbo5uyZZLCPNP
zoInktwKP+8Qm0QX88n5hvcUtIpdSYuLQmK8NasjfpYNS9tPEuq+uVJ/tWbU0L+4MMi1coC34j+A
8dqC9QO6gK2QNSZk90PWjAIB0e1VJSLZH+/p121ApkodwcLqEJAjoX4yov5GlZ4RIhH5JEqQOXPd
pG0C0nqzBnsmGw7E3QhDNh0flPHIHaJy6GBiBCM37BBoDBzeGBLMyNhvjL1pxyCPuUezYcwPmEm/
Fk/mJ+dhxWvTrT9pLehQc/RqxT4E4+3kioPk3LtFiWB7f3OGwNrHYqDeMIUnvfUBOymFPK+5bsXt
eXzVN6/B9OzfqXqCdcsZAxmDOlwotC3LVY6AVcsMlbQfo0pWgJr/GZ5EO9QFWXfsPaGjwBHitRKo
U+3U4B+zx1B1r3/H16IQswYz1Xzti9ssCIF9kOsg+PvrtoQc5/M3oOXM9Pnate914j+blzIaMEzm
Kgf/qDtbrOuktBdbdrycAYtf5bG4BBF8+xtp59BJtU+wwXb+jJe7KZTaUZRy+H9GzmCBHvodICO0
Zou4f6Pv2/nWDPZn5RJsBYDiPEBT0QYGoQzKP4L4+c2dcH8f6951IeuCNXFM7QqX3C55Alwe9wiU
6AqTyhwjtMbsy/UB8X6KpyYYGlyDD1i3Ci7UnEj21bJg27JNcwoy0LQ6Hx3Ov3tTmZ+qxqhfUpdl
DIZrveCJv3T7Ha6NdnXeWIubUssR+CggQ58Htos0wRKcb96Cb7XCk4aRCAhRJZGWctNF3fhBCZCv
fUwZ0/q3YW5fdR6mIdhPj/NdOcsx20iKunWFnS5pDKJ02ji5CHPuSLCQS9UXrL5gqxdnxopN/sz0
hnoB5/wB2aywzreB0lhHRbNff8LucQr/RE/rEcjS73BwlFqTaR0wROcbbztmt/RsQ/rEdOD3Kqp6
QVH+KOaqRXS65hVaoieSjNPuCAjs+gfOakAxpk4Y7EkvTxkZ19rlLZL5zEJaTi1gh80TXfJQrvoX
avPmxXQM9oosC06NNfqbpcl19Eh2tyziMJkBwfh2MDF6PTCrr66PdSpbQXTzbstv1g2fP/uN+iM5
uEh9GBtjPa4SuCQpHD2vxCirdhWx0dyH++NdOGOeIBxc7iM+gDiQ7Lg31EQwB5SaxtgdaJmxRe+r
fJfp8+EF7ovHfeiwBw0CwReIkIf0o/C2R4+mZDQH0EHMzzqG3bfNppfP6mimy/dN9Zoy+GAFD0H7
MeKg3QI0pkD+MxXJK1qMiTLXr+hy3ArrBdqwYdxdV2hQ3vAIPSXs2Y7GPM5VCJgMbeXMT9xsV0U5
nQVyBbItKx6K12x5WpYPukdQsfN5Us/PcCk91r2g3d+fkYwbdAEQmRjEt8w0dLWFHWDnl7g/mnI3
luQIpY5OMF0gO9YgNvAfTTNfuS/v8OfySPyb3D5y7g6jlbGQTkhr+Baubb58C7ZeGLg5Vy5SrxUq
U7IHpQmgKiAek4QGLZWATSqLnlF3lzqq1p251mIqI7EhJOa6z/tThfwowUnsUPbbclzgtnvVl6Pv
K6GSvym+oygoEz3fqVcTDPC3VMY/hwRAR8qw0rWCR001tSzRO6nEr1ZuCw/3HNr1Z8rg11ZRbbse
oCNMYmDVMv7dz86ZmjSlRJ1NReq+uFdcbYKsS9+LsERcyOTk+wXzBmv9sorww2n2izKdeusfwYWu
Z1Ksp+iIsHYNAjeFumL5vomPGfNhq54AETTPoGzNi9/Gqb9ywaR6Yl3MGWqfA/2jpOynlnh0fjYX
PoPCE6dzJCseGLhlHjWHtRhiBkZaDp0BW2fKXJvmrZvrP55BRLrr+6genZhDFxdysdpTP9k46sSY
m7ahr3cEAoDf01NY7A/TuNbfiIill5lzk1YzRUuyCtCDfhtEMuLyf+DUVG8nMP0YD6yypSXdRRRr
QLTHpvjkJ/kqZRngF3yfcyv4/RvL5a+ZnWjYquPFwgPavBKOHtV6XldVFxwK8tIk3ZgaX0eWZEbh
DtF7QiIfv0JbJJzLoBIdeuA7Y9w1AbNMw6KB7FNezGgZFYyegMM2clGaInwwk1IBNjEogh4h7xJL
yU1uDFPwqEFS7hLanNBq5zV6728HN7bj4RYLcAi2T2NC4+ShDrQ/tduHx6Juktf6up3Nz5Pkrdzn
1i6gAJ2H03E2aAxLezAztulpK9NN2eEQLS9AeBHIog8W8pSXNjPcCD4ysw3AQrwP8tuwPdXrXS03
oVAJe3dPzzclBWrLq8Cyp9Hnkt0ISmfdwNNNKkk77LvEpQt+ECGTmDCEWSZ5iZtAL6Wgg+tRO3K7
ZtYABh6dGkczEuZ5PTAWSibB+fgOlQeCiVAegESwDgPz27XpxwtC8WiC7LfP14qHQwQ6b7u2uQSS
3LYA5l2YAGF13U//LQIi6N4iDyKHKu1FZHw9fkgTXQJC7Qfq2DsQmMrZXtHK2kDgz1HhB3c7WmAU
Vip/tINtaTLsqanP6OtIP9SSfR16DYJWebFNcwutfD51KizzFsGRSFmulxWNiS45/64WpE8HcwVj
BvDIUU3YzGKoDa4aa5Oxf45OCHLS+rFTgViJMd98kkTVur6lg1VazezryKe/jTa4VyzERHL0OeEG
2XBh1ZNiexnLKmlfGw9f+/4tYy3f4Y1huU7fORRfioWRhICCaItzk8ONdwWseaZoQHcsz8cz2heP
CNBREglJDLJJ1/T5+wqIii0cjbNJ8IANAYgwdeTwTrJOz7EvK5vKYYFeJed3kI4RYCxCyqdP73sb
anj8ZBHTEx32WYi53LRwzSuwE9BFTfVkc6hpLYdtO+8Nm0+7lLd4dt8HTSxiFPL2EQMHEcT5IcoH
q2C5067KijLPukeOXUDo5AgWp3N7pNfxhcnGDLIb9agLt3ZrKeUGD+Q/bPXJsIXAP0ekEP5osLy1
/d3A45x63fmtwkI4BPalw352HP/IbRFb6mN4iSnF1JbkzmNHtlUh3F+r/LeuiZqk2Tg+knz4+Jb7
lsh4AkCoZvOH0OToX8ZluiN5z/CR7lVs0PYykgPPmQhpxudBL97eEMad66OkZgKNWBbsmAAbNUc2
/YDnkGYQPj2bZEROFyFiCtHomeuY6OAAtC3latH98mEaK9R3/GuIB5VgDo59xcTfaHzJxbDgq1OD
Ikhl3FSLiJeaSTlzblq1ai64nfuLcc+hpE4sI85XuqlwmQy/BcaOl4uyxJ8yWR7BLiZt0Ye/UJ+w
4ArBe+2cN2d8Ag/rF6wJZttRPdeZClrxJRO+9BePaiFldURgfYoI6jllYZYhUBc6XLLT+PwyGO4j
X7TQT2j42jy0qR3FfuZ5r2N5oLxjYCi5AhGfgP2S+TgnbV7qFs9DuUFeRzqIFE3Lfwfdxo5VIxLV
m7ZwJ/hbSuRmz0UgE9S9uHbjz8uO6gKWhdY+H/gD1w++kelLmZcRyJ/f78eSQmBUu02BmgHintd1
c7hDd+6iYgMLBPCJb8XjAyEJ3i9GhWP7xSRhOxs3y+XWJrzPsSluZbp3gmPIodUWejjIVZt3F8mL
dXkNGo5YJc2hBa014MRYQZ/QN6NJcjosRAq4NkBHew/Rad4ZVj9nCOAxXZRdU78YhCM5mvqj9Y2a
ialMtpdJDm9XvVZn0WaUyyTrDy/WsEws8AaHlqR7FhY3DHgn/Ct4Y0j4C52g/sB7dbnviTqXfqcn
XcLIZnmYR6Ymko5PNPyRnn+f2gqlvAgOt4/z2bw9+sWTtcCk7mDLNVaL4+6t5lyu0QmiAk5IsHUK
G/jWMu5s7RHjdPKRfrHUMVN/odIP+jiVdXTiGQW0FmhkCOxeMTnSbHS2dsh9DPYobghMBTPF151Q
bwDen4wG5F5vT5SncejeZwAAx10+yJfGeCWIoN0mzMZRgWnl0k9HbSCeCwy/Aehhe0zW2F5WnTpL
3jNLKcImQUe0wcK7h2GCcaj7oYpLIESUWlGXtydlksyae+YXxQYY7SdujFESkWhiDagOE+WnvAJP
ceuJUIbWHHizvVWB+iZD5dvVX81YZElSaz1dAzg8OtQ3P/ruiBLJrvrazo3Lnrs7tQEFeuZ0ylEq
d1HCx4fJEZX6Znzuapl4EnpoY2E5ECiCK5+TSUycRRYO4IqFPRGdaFZlCCLqieaCQ8dqdJh/dii+
1tpLsWcoc+a/0RJfAHrYii2Y4LRGhTGHIg1dDzPfkBOS56FLiiEHHm5/Rqbd1xiWQOsdo8z6s0gD
z3auBwni8qTlBxYwU3qoxtwWTNLrqUlwiKXbbETfqAV9qBMK4bwMsCaxltPwfrRjLQF9Vp0KtrwR
MtnIdxQAJbd50A+xljNLZdbDO+YiKlgCULKIGHeGZSZqOMJxcBXYbPr9RNcVGM0un589cWDlLJwt
dneLDAHxQI1vntI9r8CuL05rE6N2mBAAb6ziSwnvJ2/btrK0TTdV6Q0An/TNGmLlTyuiV8sNc1EQ
/t6W7/WUbC4ebGWNZehooR88R2PX6z0zd3ELJSDPQRNbQb5CQnaUcH0MuFy3bpEdw35XoVE5bUph
o/IpVlDfKGoMw0bylAu3OHoQ8CaHcYazBTCEXyCaY3XKglSEUO3uAM256f0KDLLl/cL5j8GhI/+c
9F3f47yfVYZxuUcbEhSwwKhr5muuJxv9s16jbYEc+A5Daqtx4EmPym4i6+pO4eJ8efHk54KRoZFG
s5m6Js18DIlRgrXKuWhWlOk/Jp0jsqF8oZ5iFh1QY017A4ZkQI8TBV9F5az+9lePl//HMWGA6bc9
Hk5HCnaQzezxpcdc4vok5//LWLoaWebMedeq9BLowMEfhN9yflZokpYlUzQx+NN3tG0QxCGhupEv
KJ/z9hB1FNd5aK5un6gLbQX0Rx8qs9AOa+Qi1cXXi2iTR27JvxtegRsaTZToGmVD2a0QNGwXKNWX
PLJ8xgrEGz32i4yUpOHzxFp+C25Wd6i3oUoSEyejj6q/tW6wWP7VBRz13LQJTjfFWvIZhP7+W0FX
O7iXqx6Q3iOJKjZt6LRBIzL4vG42BQYeEII+oznxzNxQF6+E7K2JePWNMTp6R1UgrLq0qzdcm5Q9
ytyemU1vMdCSh0v6AAbQyptWcCmtJ88MAX7d8dEUjKbvlaZFmCPK5iiAwV36lgZ9t5s+CBAGX4uw
cJvHFa3SJ1jfUVei8nlHV+ZhIo6TTZV5MT0NA+xA7zuvHo2uCKoeMLDXXhQY6lctgQ3rRyzG6rWc
qgiv9mV57PHQ0rWYMcaEWS4yYsJREKGSLBsyIfLwQvA8cFdGyyv1FltTs4+LCZiQF2c0/Nuj6He2
AVRb/be7m1dr1UOm+oWyb1/hXWFVZVFFs4poSfIDGrJqMqEOyjh6dhJ+otNMu3wpYh6QA7Y827DL
a70eCbx6N+t4djSj6QnlkMIrjdjCodVkwpM+SDoTnYYR7plInpVW8OTZVaWutdFqq9XeEaPGAFoS
M/MxM4AEwwhwVmmwwi01Zrn31pzkhfg8/8mzhdmTDYFSH/6cBoaUOkQpjqGSQcLR5+I5s1++owkV
/ChS/3UdEN9MeZcLaWD/EGT+djhQ8bPdaZyAkdFJbtY3kJ/ffmgozZaXzVMAJeClrJ1H8dDfn8PD
WeJqVwzEe9jHIiugtt3EEfTlW2j0Fa6VGfSrfcFzRh6VZ6U0bX5mgBlpz+08MOoYEqJkFJRu4NJs
IT5fPDD4hZanuVLJ/Z4V0Hl5eka+4RdKYDh/86Cb/bfB5Rl0W6We2bB6xtGMnhPb1VXMe9jttKDw
bOkEWPKp/QWkLIlqBdQCCJOP61ogaWYSR7rLbkJ4YucAMcaGG9A5CddaWgDBiJl6jxyQngO46sDM
scDd/cTqL6kh0Tbya/SXhpeTUzfMJ8gwbir3MQGq6OsOizCiMcL0voIIRLzKUgPF6AlmhWhoB+13
m+7f94JbQPI5K9p+dT9bBjmfolbs5NyX9ZlVV3Sp26knmpkcCC+hRdJou1QID3ATbH00zmaBYfZn
nu3FCXNN3RE9o8n6o7qdTST1iYSxhR3e3Rz08t35pbev5MPNx3YcKNonCBn/acGkDQYS8c/C2wEu
DeTn8Pczs+Yrl4cJf4lRAm61ZV84Ur/O5E8JWSmYNTpIId++XrymLMy8dA5EkhEQuQD+xbj3OGv6
S/OESW74/19yinrs8mlh0tKGoPLBAW+u5JZiDu4eNoKKMX5obnuOSicqxeZbFuhtpqzwKMU3xUfg
xpOvjjKYf8o3bJPyk7DM69ZT7QVGivZTmxrfJKj9fE9QEwwuIbHf5rTd5ekB98PSynpvkZrSb9/w
7hM6Iz6IHUZ9ENp1H6kRLOpOyKnir9ExNsl/crk9D7f1qSZRHTYeyGIO7ZE+fqJI75xuWwqGnot2
qHNB3Xseiu/ExGuSr8ctyOd7DoeR+S21OxfRxPUQXbqxMWQEJe9mJls8tx6UdjuQSvODhIF2oXzN
uWTup5x00bs/IIh59pI8IU+LezT5H04ABcfwlLv2ArM0Abakh1TdynCUMWCt7Lq7HZiMr9y4l9sg
BHVL90km97VkJbEBPKrfsD2GM9SR4g3w6loMyP0qKc1kwkv8Ds0T7QlnYwX0y+1JzeJ/l/gtQtxY
B9ZJN1PEbD3EmMCF+ZKbudx5h+yxy2JFlivpbe8O8vGPnffSZRFCwmeR63ocgkSLY/BZ5aeAaw7d
6FH0D5dBLHTcYFBmIMx9FtihTv/dmnubBLTsJlFO4hqMwJLC/d2nk5yFa97RI62DG59pTW7U32MT
3t5be0cwPn7CBTO/BHXnbZ0KypHG3UGtsCQpNjE41Kv1JKUTDtKbG0N1VmlBd/vjZJpu5sneP7zF
enzPFWo1gCGn0WKe0N5B0zR/2GsskZwcNO4GJA9Ss5zuzjA06CPz+jS3JU2q+nirhEbdVsEBkKq7
elY7xRrS0ErbgluyPxtdFdlqgHvDigftelYjt/x5t1p/pKs/Hza4Ue6Gvk5M4R7mKna27zCXyRJE
op2YGGBWn8YhCMfkRl8MaHeXdBQydetICuGok1WT77TrU1oGcDbcJke/fGM9i9NeB32Ja9sSLIaA
j6WtOLivV3Aw7OfnZSkscIVgAnU3DCwyQLghFE/b3bG0+euYQjMbby5FKvfRCVPzhD9MqJFC0FFp
Qe+En5HT8WzgjpVi09W8fMHtyG2+GDEc28Uxu9hIIzVvuKaZtrqObdZws0btKN+rLPTISC9YpKCh
k4jfx1Rxlsys40RuGk/6D4op32OVnpDHy9Q9DNIsGg92521QlwRKsJiq0MN42q46luExtcMLGuOO
WyoBUcZQVSBcllJrELOexCayLldvMtabEW661EkYIboFOvaYSmACceDGhvznCAwDCcFuqWtZEFhC
KQi/dtwMUgTbOzYiIukeSbdzkIYqHMs3PkeideVW0VJ4JyfO5Rcy//jOuIFKik5GwWgGY6tIYjpo
ixWAQGedV3WR49Xev7eckGMkzwkSmNs9p8edg5/UEVukNtCepuFW49H9CKCNtz6GsBHq63nagBUJ
/snu028yFl3oH3PWWz2Wwy3KXjILmR6CQ/5YhJo5ShU354ZL+BfrytjsYEirKL8+l2EXhRBPbowD
51z7UtCHazG/V3be3Wzz1ee5Npp4/R2SiwutGBo3YPaLggzDE1cg8WAYG4KLJH4WHquwYOaOQ6gm
rUeZwAU0z3oCRBZTuxUoGklCIZmrKR1IjT6Ts9P1ZZEjVM2ITuZqFOOFMwJCJei1Vk7h6czzbeSp
/Ts0uafLLd4NVZFqZZbyVpvnSN6YRn+ecmhWYw2kzox6m4v3KdOnCq1kcG8C8EhkWviNNSMaH4+e
A0fOfMmRIIbHY7o3W/TRLRrk3/+lLqRtDxTSIKFX0jAWKvoCJxE0NlaXbRb+KgA/noQQoV0/YBmK
jp8QEZZNdcwyyK9Fm9bKu7pgr/y56YqsL5Vy2kct8vm2zVNTS6TSFACOZoCbnaG89cx6bgG8He4H
BoPTynqIYsVo9FRx3zDx2dFic1hed0/U+uRS6aTW/DJItzq4WxxEn+RljAQCS1TiCnqCtK7moHUE
2jL8UC7jRNVxJVm/Idl2TitGBRKpGNy8EfiAwbKHHgD+7QJrwDMHE7OPsXGCaWC5Qx1LGESe9kU+
gS6zfrkNxLrQXJ0jWsRPk9T6j1sqox72a2DbNDC8tuhU5Zdh8tmiF/8KzzfYaiQcDqZhjqoR8qfn
rUkKKfTJaF/x9JFXMJpUHmaOhCjVeOAhBiO/uE9ZleaEVKRrhRq4/Z+t6LNHfxhchOWehYARbIpO
+hYxSGRWBRhNOokIWmDDkj3AAFOBYEoQ8pZBxZbQ9cFzZlPghL1PTRVmGj4uUpPawm5lYuyJvXlC
7ZSD35Sl+gTupa8DiWSDc1CxRFgM7VysCPWX9pcmDb+NACPaz/KW1+gSWHQ5H20iwu+Ud7DtfbfN
XNM857wGPCqVfgwrkp3PIo6mUKZ7JQ+zS9PtFv5lpK5nvfXuyA1i7fO/3SzY4Ze1n48MZHjiFaL7
mWogpp3gMqNbH6mZfcRUE7BPHcTn1+tMzbOI+4IRIKgGA6zm4D/YEOfpdnzfcpAeVcZpZZOB1uUH
8wPfaxIi1MIoJSr5/mXqgq1i3z1dhaGKG8Cbhch3uXJIrvu4AW44YcOmCoeTTFwul42WxxvoaotI
2ViWWLDtagfr8JXidVovzQF8AtItWP2OSk9F6xSnuBgExS0EoaIxS1Efiq/3FgIuFYDuPAXUPo2R
vJgVvpJ7l4Xky1g8ueMBuvNkqrdQ8eKiqHUyfNJr7i7XFRj2TVUOK7GrPgqpTtzJpktpF0H7+qYH
Jopfwz4oLo/b22OMZej+N87sKS2Vj1OCHWNsM2V8YcXbOPeMrituu6iGegVei6CXILn76hAG819a
nCzqzqDhrGEC9d84MzLKoOgdB7TH2OV32WwHCO3JkkOt4DpJhkh39yLhCdxSxxEkF1tmjoCeYRYo
c1LHTPOppnwwaoIfJ5N6sqGE7zx6XfSdTPqCVoH0nPWypwWqXIvNU0mPqK9SUxGYjMOLBOC/6jP1
rIW7VLTs74aOjVytDnSbuMIA+Cs7Gj8lZ4i7D5uSVTjr3If0aCbnybQTwPSYUEhfr7ox79N+mVLx
C/1EZB9Wj2C5HowgVWwttcVel8zT0x9bV3NmhGrV6PKjILcNxRNtDLXjwvpOz1yubNQEjtMRJZZw
QmiCVTEuWHxAJ+eFoQEZU1R+So1pZAsg5qmhfWZ0iiUNNVjrXJ53euOoJfHX4Hte+nOTSBQ98ePN
DvWyA3uJs4ujaLuKd3ZPlU4oaaHS1/kkAE5FkUNBucbsweyIRr6YFrAY+wdmYrbk76w0kEZysZYU
73KvAM4IXO9v1RGIqfqiU6IyFnAxYuS3+BxGRY2G9jjwfi9DCczHYzNPvzEOoqac+70Dz9O4emZN
GvMgDiUbF8zzT8s76kTXyoTtJJ4mKEVPCu3slT+3qMDeM5CwueAF7StdYJ1up9CqsS9f/ANVqZPz
J1oM8O6+6Yaep04CQpMvTMTwWOBRsjC2I7Br2S9MzvZHlOrh+YmW0fMJPkBp/Y6Vwu1e4HhHwmfC
Jgbq0NWQie6KDno10c1VzMfWCaVigQNOVmgwmVz30bruEdEE9lHObLIOx1iW2SWFi0mmdty7ar39
m0w5p3wrboL/gXtTForG/T4Z69KRzfyUCvtuxRt1pIivdbOYjkIRDtylub+iNF5uWNNehrMtckwa
XTA6hG8NgSFZ6Lg1rEnNUO7OyaWfTT4lvUJAbM0/BGQD1VcyXkMQrVdI7tl9ULWLHXOhnGHk5u17
u6CifQzkvwWREaRdOnFC+L8DHKp+EvvHz4vQjTICkyLZ/vdRhu2JJ/6uk22KuQ8dsn0rrN3SWonX
BcWrMASI99/QE0dGtqm0l99ZJbEmPuMnqMvTzFIKhxGonSpuvXfQnXWwj0B6Gr+dv2SeDeRQoeMI
eltr5ecrBtQvHDxT9JQq5sxFRnbg7aNg7J6vJpe+2u1NLn+sKvg5ZJcL6awAEEN6rXY3EOyRmh79
ZllQPmVPvShVKRC5QCQVjNGw2L4Uq4/tC/r7idD0CA1xk8ZupKcdNN6voY3IVzUdEbEejnpoBf3X
73OAc10xNYkiTWhUsRkfNPLfVakquCmpdn5wRvE2Sh9WmOh6hWHUv0AagbeoP0WACLUfTRLVwn4H
t6b/2qPij2DM+VBaFNdBabIFzYbiZIJRiPdYzjphVuZWpAzUIYQMuJZUQFOhVzVF+HdKrrMG+vl+
7RvmcrdoaGh+Ji2v68Ouoy4Y2WYkm265AMMoZZOVY05zm8Toficd7x1XPmoUervtnIrTpXK2X94o
ypbaPwHBwbgAISSU7T6k9CjcWk7ga9mcM0tVOpbApBjXFRU36FcLRtDzny77QL3rG1ZhmLTkY2tg
OqOeiDK1GB/I18tETz/Fplh8QzQEZrG4R3DODAz2VlyqpKJ3pGzddWFNI+CDCFD5ilOtrp7Aox8D
iuM2dVmHklL5xh/3rsro86bn4nty+fVDewkwXSghXlflAm2U0Oa+ndGDiZCkwl8lBsCSK+Gv6tTe
0OUDGf8X1+Zfst5NeW66SliFj2Cxle0skRkU+RUCnsfSEnKS1ABi/R6rN1609PyIE81381JgUe+O
ZSo2kpZIab/Fr8z2Nn7RSsPWRgqa51/rz6lCW8DWR33TgpnHXVZBaXZGEzQ8dhVDfkZDT4qlGjLH
La2VDrwoOqe+DsST2aWpXOFJhv3oAY9uPXxyE6Q/QFs/zgideYJiUdRcPhI/2gwxIVUytb63w1hy
p6SJN9uy2+5AQnIwCmtVSN21f7ARA4t5iYMF5IWp+gTDYqYpryMqEZ0TrhCSBw4P+P6MaghLuOwO
zrsA03GORLrG1JE8hxCAi3e1tfyw1QyiaV7X4GXHtCzuPa1mykw6a6kE517mwfLvc3ejw3+4UAFc
x13npYsuHiGURtghP0UFv0jjQBSfke1QiD49XW0or/uBEvmeruy3i22nrOpMNfzVSHVgAuDysYcf
/GGSf0+WX7Zw0emz/Kuu/bQBU/xE4km4qOYa1hYrrNcQG/poSwRVEajJsmGLquzEgRFqP6RQ2GlT
Aiykk1F+HDU2NlsLSYxepMhf/0bTNYkY6YpVqK94CXhTan+zKLj98hCPaA1jg9Sr//Thn9FL/lNV
eIekLhoXprGFYYSJyw7+AP7geD5bvO9mFiXcfw/qbDwfGUuos1ysvxBD6ybKbbOMDyhoGrWLnPGZ
IkeXJKHZhjAkm3S5p4envG2a5B6Y6P2rJJQDXa09BH0T3K/qtuCz0L7MIu2lnHtPqv2qn+RWptRw
PGAjHrUzjFtC4W7mCLmY0vXkBF/eyprNkKtH1dvAvnyun5ACgJ6Su94UiZjt5dLT6BLPAvc+Bmit
rUfMG26uCebC74sVnlHDwYjJ5caYAmetyhUzD/bkZkEiQS8kWYmvHC0+ojeF5FRpqcAe5/M90DIO
qBckk4ua/Ai8flE0FtZR/3Tp6CjXhBvgkvYmvWhh1Me3HBcmG77qlb6n1LTCOtQ3RStwnQ+u4AGK
ub3cdtA2COqw09vxfoJtJwTdF2YKjyNQWlF6LGzFuI14iErhgWRnQ1/M3OHOnnVrr6aVIiUL3Okw
0BGc7AsDnvxu7A2tpLYArwgh7Ha9nSezcLndvxUrqQFx+pV45k33BhzTLq/6vMVcmkDhwdEtyjgG
OGTCj9LWC7hy06/c4P6EshCgvEr6Ssy8aaQT7Tah3FkDkAWTxTYUh8TJc275PToiVE8hHisHncTz
ebk45EH9ijHY62CSzLVPIw+VHSWAvliQMK+SaUshhTS8vIqLXLnzDMFKNVYCo5uN7sDlBnA8OrEY
OMpF3chh+V/bJ1i5JW3uTe+wy1owcOR1PHV8fFUXw/gu3t0eu1PYOAK3pdgHfo+cGMU9e7D5dgwk
F5xEyTn1Tf3HzLMyfdNBo6Pn7ePZpV6UInIVcmHyrfnmIiZwNLR4iqfMePVuFVGoEiJYqRfCgkeI
7Yh5QOgsnR/zFe4SaoH4j06K4wL/x9XpdiYj12hTPpx3+4+kyDNmsHZdl/Z2QwQu1Su5s34IPOTs
hMQR93+gORfzSXIXQUlJEuW9mGR02HlP/RPaXuWlUIuRs6l9r5KOYEe+3zqHSauWL4M1oumtL7sw
Vl93Z6Z1mqQcktvmjNZD0+3AZ7Wgs6pp9t3k+z6QgRPzOwYWMB6n+/RINXsEG9pHN80rDcaeV4Mq
6GpLikq7GuJVVJIlAd8gNJm6R7WPGJZdcGUtF/dUr30OE0ViGAP8tiDv1ajrZMkYvGawJ5F5Deef
xKMAh124kwgz2Fv64LiUarYUfgnwv3uHKYNH3YVrCPy1Ar2OOZ2rfMWS8H+Ky7LSuowkkFW3YO25
35lxdSOF2ha7oED7xEW/opZgzqpUIOg4wORt5+MRSqFrdH1eOaDpw4PruycpJeZ/3x7bqAV43FFH
uJp0S9rAc3cGprwB3cP1fbGv7UYIqdEb7if4ewE8CPDMkdllMjAeMkJF0JcQ67pavHRdL9xIizlX
0QHyR5sJIeBQ6/7T5+ZDeZPV0tiwUOoX/p7WyUc8sEHpBJjHfjIuv1cc/QytB9h4XIddjE3wV9JP
JPX1R74mZYneAVCH77V/KSXrDqw3KLdilbRtYnFZNGAi0N3Dhlo4VlfDV/fVik+fnCQ/Vqs4FnZ3
AnCbQDPRaYU8M8DjWGfE5jXAh2iY/RStuQuR87zmnt15x2PEmwVLNRx+rtgn6xyO8LHFLTifzMGl
CoUg4WORIAse8jqKXaFowyZOtGm8t+bmj1/apjwm/YF4nNTg6oPoFtSF+GyoG9Q7Ui+TM03d1/GU
gfrK/sCceJ3q7M4OtAOPLP1tXdpkk1XEybArvSAP+8Dw+fcOmaubeQHqYxVsDTibxzmCLcmZ+zUJ
5qHu8uE7LKiQeLDPC++r6usYfdI3aPYv7AzZ+07GiK1c0kdNpfcwW+hc562UNrKmb82jSYecTis1
CwskLx0wKivxs8coVr7VvmaoKbLDq6ZM2ufFu6qt+2mG4F7vewUf2caf7gy7Tm56lG6stEae0plk
SWtEqfnXPgxMqjbyZ09rXEZxoJuM5NDVtKVXOCbCDFrAwFvKB788Y6Wo4zAyfRSQ+8HBycewO4yR
tvN6V9NGvalyDLytc/VYK08JUNBbYDgSwfJ34KnQOy2Vh5YCAfjDXP0RWlwXQstkgejXeLvkCVU3
gDZclCpo2wxm0ejax4PiuGv6huKV3VFWsFUnO7iBgKi/s9iHirV8T3MXams9equpDY1VI1lYiIZW
n5cc8Z/oc8+0/CiLG4rqJ6UbDUZXI95f57NVHINNZs4MriqSkHalxgVfjHdO3CXQXNiY9w+I49YX
/JjV92SrLzvmI2HirHDvgP9FTBbGXsh+Y+ZduQqxgCxJwwKY+S1ZkzVQ5+HifUcV0qh9m/P6GaiF
r70l5jSmLYUhYsbsxPZZ/bcxjCRch5Y44G8K4jMxT9U8W0OjPfloGoCBqxHkflbwhySfqCdHKDLD
QzpykJjJmjKoMqpdogsyV4luDQu9gTLLG5y6Dceir7iibmvvygv4MUqvnNqGVDWzxpHbjsgnK+JO
yKIZm0w2zWg94Lln4PCGgfLlbQO0ryzinF93rlv/v7qSYCsgXygMtTZmBw9Il2eXVJSW3JCq1Mb7
YeXL49lR6rHBv8rHDDCfro1BK0++DBxowADW01kup03dt7wV9bNt/q90ysXLwklThmQFMZxmdOSn
cs8lI93lHjm1Lw1C+MKYlW8xqlHGTT3p7MUHKjrrWZtdRNcRmE2E0ILPmK80Bhk9j4aUcXK0iv3O
EvKhc26iRuecSu0TPupU/Lp+5P5bEQShLFL2Aa88YQ5fkZlQSWXox3doHaN8FlPbvZ3bM4Es06lF
nIqt6QQjbOdSz46d9DBXfVq9JszdusWU5/3xoQDTS1sQNNl8OUpaA64KTAQwikk9m4tTkS9pej1y
QE8hRRVSgN7EBGa8E9w/K/HLiY0xD4K7fiIwddzWldSvw3VD1yfzzF6Ni54JRINt4QcAc3DWaL4I
ABR5GfswMdmpSzlQkM+BUP+4mBeY2e579km5HaJCIucj8wsQNqFAasyKbHGxnqV1B2A2JH2I+dX0
m6viICqiPMJBvDRokEUIX0WRZB61BxFU8w9uSI16N/EistlkvsjcO9KYJBKBpv/kTwy4BENtxq/8
17LheOHwy31XNY3xboIyhhz4xp0LCSVn8/+t5TP5V3faU4x8lUsWeEx7rLhUKx8bOB7O+cGigPa7
YNA4gSIe0/HCvHdT5A+6PLDRY3tnRyC62JMaFzzotvYZhL5GDov9WqditBHJXHoU6jNGK4/yzTeI
doEWy0y8Dp50Ofni4kxoKC0PNAaj7UPsyqvVPgyy5z/UYwoacTKOQafJqgb2R3DRZGyiAOrjRNEF
gtOK6pcY8C8tM4AcXUn59PI3zCWukFvKI+dFzVrkKXDwd/uNaf2mUv0RhC0Rgxy3mp+8Mb8QrJK6
nVAKeIMcm58eOJEth9r6tkbF6Hdkr2EYwX5A73H+tta3uaY5laoWOAqf0lK7VomJipSnHOmQZvUJ
fYMDCBojs8tvxRIPRCKyOUn9e4CeWY2+ynZuyrlN4z9t8r/TgH1+ckssU1R/uzBzjkMlXGJE9Fg9
Etju5fNk0h9Mo/yr8+vwXnGM5VvbJsN9iPrHjjct/kBKrjx1v9UwsIjAZ44KL4F1DxaBemETqMd9
o8NlixcABnhSHfmAPfTkAbTgHwmSpvXrQOKPhlhss7q9m6kPJB9fIHSMVlnpgsHYTVBVUsiyamWw
U00jZW/5iy9mEbX5IRBwMMV4NcVRxOZTyHopK55h6WjWdCQZkIC3Cyl/9LclKTTn7z5kNNom9wya
9bratRpgoLwhabtFuQW43GkKUnpeWYTotQYjqAIL/ibaHyiywzNh0oe3LLYNCtLc1KK7SoBhCJ60
g4va9W66RQM6qKecREeJ9DxeZvX1bHhXOLGxIoX5wSx3xZ69g3P/mAUsVp48LUt1S9SwwkFYV1tr
TgCKDIspj+9EL+Cu5g+bjyUw1uqEs/xeQ6gxEJq+Cfh981su2zqfd16EDe2lKbPIwdEztkSeFUKL
mCWv3LsyJmRLWCljUiSjOGgv/ATHbjGIZaaagFHHxtdZTRo4sS5KIc5wDgQqqC+3/NNwyJ9ebz+Q
Y/QaO4ZzU0dwluJzdjC2u5uhYrmuF0hgy/HV9J73HArPxz9+bWcTXzOt2lg1+3gTNOoDkI5HGgB2
zVl0mLcK+bT+jBDBjo0E89dyww20ay/ba8dfUifgvq4rYcnwsB0OXn6ljh/uayzE4M/vHjR1VFiU
WU8/9j+JnHf5gZPmU4ne2CNM2Cr9VRGa1rpK5N/2DXFJnGPD1gRLqucQns5olGIg7MN+knyJsEJ8
qtmfJ8tCTVZx5F7vqZkhV0BuAGbDI3+2fFAw/bwcbIF4fBoRPZbU3ClyGVZ/nOSXLJgMBZ+ZXjW9
48uO05Ow+YQGDfIM8FIQSm/Z2b7ca2YuzkfnXMSytEDACkiyEtPZJeWzBLQsqMxV5nlOw8LfKHYz
egGdAyOoTdcli8SnjVisbNTSxGax0T2DJb3IS2dxVX9RO+y/5OnoWp61f3+64DcCPSZ1oijNxWU3
MxYSr9LWr2Dk/d4Ec6gbzbrj0AtWz4gpTDarmUMrfEvtASIL8zubgvY5IM4Bpd0XDWZYXhiwV2zc
bsP65yuwB+vfj3ZxNRmvUYWsxobIohstW3gTyMtlB/C/x2xYk4MNWYlkAewW4jH8g/DUaXHz4IaZ
RQnx3yoNrHU7yiXfldL94h0TgoDz2Mqdowh0KAu7hdsuQdEKzNCtf9j4+lBlSpmelkEycoJoNVTT
NUAqH+kdBU+M6VSvayLHY90Jcop34zi46RzYg9ZJ9TBblu9sDCOet6ccgRqI8EHrhFjXEK33ALwI
URJ8OdmrmK43Wrq1N3mpx591ytATyLHf28+iQguafzZqa9KnpQ3tLEsyAVW3amQHHwiu/X4pQ0QU
bEucX7ewvbuFaDYvIk7ZJ1ehL0gfxy7MS444XmQIA73Nd08Q/q1N5kbd5LWKXFdTbK0MuRcngrZt
uwSulyRsu/J4mR5uNu0Mxjc/gBDDD7SJ8IeQxXdaFU1Ejlw2VbKqREmaguhnKtYsXoyhjSSas75D
DR3LD94Pzw2LetuEqTCSS6Zq5nZxbNmDvwANiSO32GoBcojVCDTcclmjRVxamriHXfNSSuFtF+1V
TcHJ84Lf1Zhpg58wswWfjeZzGbmKCwA6BKK3clWAS91soB6p7XNl6O//e4UFiQsWOdMEYHghtw4p
oX0hjh4cPsCAtobFxbw+LryIxLedpBq1UA8WlUeUqxv2kz8YDwIIJXwrWchaamEDfYYg2c3QGUi6
rFyrYBw9iyMcpulmAeiT1Z+MmkDkD28vSAqOdc2h0FnjF5k5ix6Vl5dtEPCZp6S9Soms2V/x7k7k
JNUCFXpkJ9h4qvwISUGzm8Sx0G+Om/O1qJ7dbn2aZ1flfUijD4gpg8z+kXy1Twovzu4RyxKw6spg
JyBR1bLMkYq9+E/vChWk4uCgJb9BASsrhi+hKlgXxSyBPDKBbmg59MOxZyimrxlAu1QtiDa5gQBU
QWGy7bUJ0be3mwNG8PmYpr0qLTJEnL5u5JtsTwI+sIIymar15gsuR1LonKYYzAEsl0mTFKOywrPw
XGl4Yj+7bCjjO6ccrGWYV40yTSpKflMrPhs30rzAKmrYYxZ0xHNEhyY7Btdn0RBICi6vk+ki/Lap
P4vQn4n3DVn3eUeuy5FBE96xG5NKID0Y3jm4irxK33eYCHsagSYP4BwJB2dIT47FBhtG6pUHHzYT
hrPIaoCxlfGTEWwMuBp11AWwAqD0R4sz2EnkD1AA9/b3YEzagjKG3XrdQWGILKvJhRlGG2zsbTLt
dBFHutNmb1pOb1DMUckTHxZw5WR0XyJ600Y7sUIKuRBfrSzHBJsBBDF3cIdR3onYTl9H5edX/5YY
2ruOQTQAaMh/K7i3CEYty+3oCJE7DXKky4R4HhkfMn4ANdEvjzdszRrMX8KgF6w+bA+5JCpatJKI
hByJGpJNE3tRTxJcHdfePLGXNlKmN5RiHXL/oz9zNZvEfgT6tapoG1n3kvCWqe87HMct1lvkIkQq
enpce37u/wgj6rqXaeert3kvIC5hWkueIq/fONs24nDqJoLcEJ6dTxqb/LEPHn759ZmfqCLIzIGS
/yKRohAPnHHSfUVIH4+J8oc06j+XHSQQR8j+T0Mg60MHsxH0LNFN7vu31nBhoot+N9yi6/Wk3m1C
BaLQ0Ln0A6yPs3577IO3TVXSNn5LaUiHwoQf9zhhgchTD1Qc6eVUwNKm+vwuh8xM1q5N/4mMDswM
rUebk0jH/sk6uSX4248OkPIqDCGl7hDXrrOSHYaQPggocDLJ6bAJ1Ncu3FRLAzNfs/VvjrzyGo/B
IGbyZfK5Ihqz1d1M9q5mcbV73DdebORDrROX67Zs7+75MweG+Dgc3lpL3XJKOkf8Uyae/I89u4jq
DRTQ9SZ8e+K0nbPCgOcOT6kP/oft4xVGRtc6ZKupj4oYp+VJctIEXFcVmFR79sr92/IiX/BIdZfo
OzblfrzWJB87VJ3BKxbc+w6lRFscWyZxGKCvBcob0pSooS9kbMfZ69LuxHtYvBeOKhgCYB3cvhiG
YkVeaEm97FyPPWGwovTxp5oEaFmA36eFfF7HbjVVgKumq7XL3+46DUJfmnc0wdEQiLPPoPZGrMeh
6M9/HbkYlfp8hdyX4TlUROGIQ0BzvT6Xspn1UWulY0sz3lso+W6NQHM8Aq3BqmZZ8ewfU2Khuev9
+5FKZQ4iyNrJRzTQA9SE2oDGqGcqTtx9Wka+ZasHKFkzOCg8sdUJso+YTEAeCfDTxdWOAyhdoZXr
HfNvSAXdsVHbuuqLfqi5ACuL7sWwBc6jiUzJJIy4A9yxvrep9aLTg2rV1CueW6QvOh6WrUvb3pp8
fzYzKSpPy3oLS5PXCq6EzhpX3gnDUksejG2LfjzgeA/u4IYnXno+UI0NypMptpCFJXujUhtr0COc
e8COl7LZrm1+3L/I+cK4GinDmNNwMYDWfTT7B8cNuJGlxC2lVEz8frN+szSNjqYHKsklv54c3hLK
XawWBiDh4vjO6Ml262PBJ2NRGE2cgEBwqnEPME4ie09X7iTdPen4JAPtsa4VwgZwIyX3pfbR4RiT
NZ+Wq/3Ywy1DU6O0CNJXpkOvbVY4sG8w012sYreys9xYk58qXA2WM+KDjRE72AUy/3dROZihzMPN
zhYhwF2EnuSE1rRsLWC/oL/0pFvujudqfTJeWQQFCk3fDFZ4l6D7wN0K+48I+Qf4npYWLdPbWXq7
QI/czIC574+S1WVabV6O4hakJEbI4R9I8jYbynPwL1QSdASBAtKKWfQPoucjAWwvjto1IzRsw7Nd
WUi4ywO8NrQv452JHu7+89/zmlLiHmuDwO6NJNqyo/lOa6FmNVteOBxafNxiK3Bsn+Uddo30kuKv
/svZK9iLwVkh6FErmwyLcNiXziVQku5KpwpQqnRoDHvcoOIliQCOLr+mV4r0TyqICSrbbX6DF2Hm
EtkEjVr5MRjV7Ob4R5/gHMXe3tjm+i/LHUsnnvQWNqdSY9vIwIdA/jfoZYBaOJgNlQ+qlWH1RRhs
xhaJ31s4WGt+1iHhXx9vSJyM9YzGMtHC/jAt+onfjLYBAevJLonT2ZJ2pfpWpQHPyVobqGomX72u
M3GZoFdVshXexUIR61+rxxDsV9V1r3Dtc6/CJrie1BdxMnknoJVap4EFHHzbrNX8X2r72ScBYzOo
IEcMmuoBX2yqVaVJGZulHQ6MhrkyRJN3CBksW6P+N8TCuBtxDmJ4NuBaRamdwE3d9fSn4O6JLEv4
4iH8RhzvztC3vkTf/aKRl97Z9+zoDJ6JKKMg6/EqVvUu3rAEWhluPFct9bFuueY7591KIz8MV3Ar
INBjykCiAtZy9mywoyKXo8lYu1X5JLEA1tsMHpIpg6fOwysoeXE6tqZpWsL4+XYX0LOBAiLvSaIC
fVTc4ffzWgEfdL8QtfDyV++6sgKtKGMaRa5XEQDoOV10+6MOhwmS/KEoNq60QHVSuNh66Jb1Zf6A
uQ1OnxyFmQ2b3NzE93a8WlgQ+hxXwDZ9ydp86awRr9/QWCst/c/dyUbY8ZMqho5EbP5V/vNtpOms
47dekmie0IQ8mVydmrhHQvyw7sZMKPsAGOXLCnWI/4noKmTaRB/WBwQvXPW2J9aLiSUNMhCLB2/H
oNxOaQwM4QPQ53/Of31BqXI1EaqQzaT7svb7jOgwZg9BXV5osHSAXopyyQQCOt9whkuNlJG1BNYX
lx/IiB6hQlRKrwlD9byA8YO40hwuUAqxm46lF/bcxH8LOP8K7O5XO7+79IDEbE0ZXSbxxMZQ5p5C
4DjpOELcP9YXiZ0CCCkAD7NoRdie34JFP4RnMYTULPdMiwRLQJHYlGfxDFQW4avky+HB+tVBtAgu
asJX8an1tj/WniOoCAn9PQnxLrpDH0y8bB3Fzd0xFxTaYlMsF/RN39qryWycGE5nMwwsEHyhlfM+
eb/DjXwOJ2umbv9lJ/Uh16nm00zikx+JES0LFu8eg9K5dS3krkAigCZFMUJ1fRYyYvu4TaWL8S1v
D9GMxzqxNdp1bHE0PbE7XR5ygZNSQgAbBYfjR+tqBPgT73krdSVgCZ900t/jaZWWwz/k8WzLL8nV
rmhpya9+Z904XnAqidzwYXrZgWBK2gtE85zkZ2bjt4gdkWwcDUT5WZDntgCK/1h7A6tbtPVwFMmV
bgNsSpvF9XKfabkKj1R2AbhuTMGVOQ93SPgZg7v8g1CBwlyGrYcvtCs6tehxYigs4i/JSyStPNVy
5StzWnypyoFoeg8Q86RK5NatIjBVlkmOZIKOl+NGBnoaFcZXn4v8cF22HQl/8U37+PkwKSyyen62
eUPmPuHJduR3J0dro/4gLXjb7hfqQ31UgvadbfFgTy/v/x4bGAK9eKbbSDaksV4Dp+GEqoh0vr7D
rfw2wgua0V2E1NSZNmlldPZySJm032+ByjnV1pw/xDkZHZ7WEslRBny/RpjwmeAMo7Ws/D+P6kKu
x1FEnpwfGNZaoTQyH3h2oKu1zW5+sToD76iHtKd/gE2vTZKp8D3I+0six7Id38dJdNWKb8+8lQfv
XxXffl9gtpMoafwHgNJ2QvO5lQ238jQegANphoi76XqpKLRE1SZaWVIoPPWDc5SnA2FIrhKJVAZd
hAy7jlLKu61L0zVt64A9bOz/SH8AiG1e+p7ECJCmI2wiztJuNiI98iOS75tCZVBqc6CITCWgYgMM
eJnaS0ED99JUH1HzUowGH/mb5uEmXD+wvHRMdbuQZuNI5u8FheZShEMKYvPoqzT6ow6gL3y4XJ6i
AQOei+7O55jn9q2pFWNSxlZRW0FX0UaqHccNAu5Yj7oCerazPPcGFny0dgGYHrOyvmgPMG/gUwL3
BE+G0izF8xdHwdkZECzvDUl++qB8GnWRmAlPtxE0WemwiJaWAXDrYjblWcg8akTle0FiOyjJ1Nrx
YhdD5sZ6HfMa1/D/GlCx5fdLFlHfYNf0iGZye+b5Jt/l9LjKN0rWPxRKEhrdLYST9eRto/jr/7pr
83+4CBEyc3NumdkJOc+0i1ttLYGaPwjbsd7XxRKWKqAFWiXxKFa80yp+Z1WbJ1iDcQonNBh4tyTF
URYT/iTKmDQ9o/8UnbklVYxNamisTXXe7rmVvzg7t1N34gR7Rb5DE/jkWrY/0Qnt3xEaQwfxUEsK
mLMUKN7a0KKrOHaAzO+Pv0dWVJEFDANP8+e1VIrEm7qdL3c/LEA5szvQnBvcjADix2SkKD3Jv5ba
PqN2DAddn3HzG7dIpbO2xoR7XYjAfrXPW0Rc6/tulHjFqMKhVnaJhlqwJcqUk784119ZjZUPA1yV
V+REWb+E4jEjK2GA3v/eYBxcMwZnNibDZT3sq3gj9Cj9WdSdPiUPJ4DQE1yQNSazB4MSjMBeheYH
amln6pqyoyXh4USgdN46zGo07nGH/UQZSr4GcZ90PDVDPtDLpPxdrqVIQYJnmeUFdY+frbbwv6rE
Mqd2+uPx8PyWZ7/KMVZlsFIxSyURk/I4VNcDzjcnm+KK9OU2OPGtcZT1lkD836ZYG2bFVVfxxAFD
ToWTVqOSD1D4jT7ZpADByPV52iMRhC6LyxAky7dcrzkoxdkHleh/VqA6UXk9UvKfdvCTq6PzKw18
A8aLzwjFimHEfdsY3XlJdw9pQdLrlBo92KR3sw/YSz09b3fco4CXHJDbAAqjfKc0/sWJeUV8/OcX
ApJZAQA3/BKkA/lg2llnHEqEpWLTJhZ6E41Mb8pl/YOV7iUJCqtuoBZAHQgGUMERTF90SlcwSXyD
Kw2sGzaQFNCX++nMjFT4o6CK5ODTz2u2tEXudGq/YDkA0Z2PvBamq2FgyOGCDlZPdAARvfkhxtBb
BowUMjSiELo896RbAb+hhgO6cCiiQIq2feK2qR3gE45YlYBp65Ft+P9q9Sv9sSeJ5j1bm+guu3PW
JUjJWaBE5oL57lXl2xGGJroVSbdrYQDNjtoyih+4q5OXx8V45wYS//DWkJEosvLCAc0N6X4KSo22
J81I0H+acjkVrScP+dL9sPciCXGM/1+dmnP56MQb9aYKFmNnFaNI3Nfy1iBs08YIF++n7U5hSL48
BqP5cWPvflExHWmTo73vMkap/osl/aauMpy61t8tILyl3v6LYpFTRcnYqosIZAqG6ZnTJAOCAgSJ
0DuHtKseuTbJY0o9l29Nps2+Sj9zhsywXJw9eP0tJ/toUYtmYeRrm9BIiohPbkbtUMXJZFE8qGHz
9fOb302zZljwPmmMgJbrdqajl2aElb3ZvQjixUrCxhR63ueMA5g0kWEiuglL/cSVBaLft7sLACmo
3b01Qn1+xICZ0is6g0l1m9UxFI6MmkiTnconKThjqF+hjlrrogotznVryD2/2llOe/xu30EEtuVy
MGjI8AdDkMPJhKg6sM87fpXebo/ZTE+sJ1rIxRzvdhmxSTNqhyfnXveMcG+ZRDExzW4j+nYlzlUD
suyPNGpbA14IVtCGMZ+9bLKHE4Ll/cgvESTyuD9cq3tX6T7LeuUcWmq92sm1cPgzolY88TnjJWlW
/D5RZYv7cEODatApDIgyZ0ZaNx3x9v5e6Jj2CRkZp+jKOeOE3WJ2Gd4To02t+l0IAhvo4bM3UBN9
eCBcuLviEkt0YKGLAtOF+44CGHt7m2SOuBoSoarVEhisVLPSpQg18O0/RkIlHzaE7mZGPWWt5erJ
xWuQXFkAJZXhAPC1PZb+f5F8UrEpOZv/Mql7cHoMwWYik/8YnIbRdV+pL12GtSzY9qwZfu0JZlzL
KWm3Dse8aLfBSzYeyYJnPYX8nGlMVEseYfghAYAnbAWPuFxGtV1m118EZaPYqh/7ESZgvy8Hwk6K
eL42xlkY2toSWl+u3LMwcoRi/U6HFpNIEw/dokbZLgUIEVcpICr1AheumYdowrupVurOGBZYYy6P
PMG9vG00/6DB7cE9xjC/FKlzb2dvIgquavZjXHPUEk+Cp/38RPmuEAtH4amsdsGQNFvCN/Y7m1Jw
ncQF6IhdAeTfIYFfcf1rzEW6EtqzpgNzQkcZy0VJ7elEyX9pAE10hVk481ZZGpgDrD9208Azvi/S
J395KY6w01Fp6F5tF5qT/6uRPA50ASIgKgwH8vukfztrK5xsgXXAJ5BQiB6RPPBcj5yuISqMHXcO
fltzOAsK67TIqRk7PBx63tmHIIdwEFZmA3XnJrpjPOZih5t10ExrVdOZO5SaY6fgXYbZSyLtu8Fx
avVAsikvgUtvl7Xba/sUvkX/RqboC9Km5ki6YIBhvYShkMgGQuua9ATCtqyuoBPayBDphWH/IbuA
HOtdUlf8GwCvzD2Tw1MzeZ961zvc0E3ZEcuglkWNIEFIgor40ZzUs9BlbAClU50lnAtXcz9nMO0M
mSi0V7DhKxThogYAmsM3RQpq528tGoZ4+wqb7yJLlGkuQjlAAxGYzygtBCtON+JA/BIkwXAfqhHC
JwFs85ZeRPVrF27PezRHtb0C2GpVi5VXJY0Qy1th0rCX0ou9nQieYP2mHbVw8yZeg9/4y7H5mDzd
XhbBoveS4Gc50LQx015pgJHzlOxD6pCW0cDJP3uqjFeE/iuFnaCmIcNRDE5EokZPJk56qlt51GkK
beiw4NSgItM37b6ZtAFj0LZaWXAUf7kH+6Dz0rerzjYEqtEYFq4sMm3QsIRSnXCXsB2siiBuAkMK
jp7aBqjRKQDgnu9e7V22lHs/vwwORdJJ3yoHWoIgPPPtw/YCAtIDpXkt3/FmsTbHvhJIqm5hY01a
NISYuJJC63rl0Hl7DYsZ2swqQ7uTFSScsgIVniKZEDcRaL5cMBfXU4dXRDKOcKPhlQakhhjLFtuD
BPkyQ5UYh0Jj4nfF7p2olkGCe/lRVzDoyxUqDd+SvbwXoBRE1ldO/jk/hZN9CPvDuWJJQWPLYY6x
0WMXvMqYih1JCyXMHByv20K0AFWO1M2MYbm9Fa1t2zZR6Ikk93LZaXnx949g7oe78CmGVhDONd8d
R5oTNLWFG/ReUl1LmAlz0/AQ9PMDYN4KlecTv3fV4l40OVBCzw5rrpiVe0IgPYDrciSOi1GSms0l
VzSMzMXihA4/UbiATNV2kkTGjXPoSStVa6G3LtzV2ID8W5OCREaYhbWFsHtpyJAxQzrpgKSUGvH/
Ggy3+z/jOqABrAPWawh5au7jX0nGUB33v+DBD8P5ARbRd9sz8KyMpQPYFIpPGPn5aRFiTylY7cwC
aiDfefPNnJR8dlZevNIdzK18W2wDJPBOiE+A3sZtKrKuGG0sgSmAL/wvCzwpqQtIcCxRSKFbecR6
AdfqOHtJHJmqN/9Se7j3sIM/gvucLEUbIW/E/abs+wh5OWkKvW699/v+pl6EwpCxwC/k+0/6NWPB
ocrUGLWWOpyGWvjNH/au5mJa4VYmvZQhZRbdd5OJGubGCaCmsWq9BF035F7btarWAAaQa0kWzlHW
6T830hdoVggl8c7D1t2f2YgSSfezlbjeiQfBiEswiAD4dSfVV4OGa+XhbxySCs+DZGPRNMqkSx5p
Mce8M2LhPcVKID2Bxt4FUkocI1/0V8foorgGXHMtlZwhDY8KsglZ56Lwcswg9KFWEP7q+mH7Hu4E
tGC4lkO1TK8gnbfKxr54zPgxGWoN5ZEsX63WwZLlVIqYHo3Gdz0xYfVPrx0mVL3ZE8iAB4+jH3sb
YcYGHLdcLl4iXdQ+7+0rthmu9KbiPEopB1mFxUIp25E++xNlxJXPa6l3iypS/wwNaIxg2GvWXO10
h6RFMBFBfJ95isFVXh9CZiQIkC33s7nozeaTCaHcI+UkymxwHZia3AHibbTa2bUiniwvp47seU02
TJzk3CrS9KCuzysU537SVpDrv9bwfNKkEdSI2yBFa5AtNP1055AV/aStKjcbJOx0Om40qpPADR98
OLcCUikL3NWX2wJYTfeLn+Ng3PSD6InQLplsj+jYbMFAEn0Lm0v01WRvOwxwdpNBzMUTh/RJgWz0
GdU7mFp8zcqT02PGshE+GpWcvDgy+JhAscndzKAWOX234Mq6NiXrDOeZtpx+8IW4CI77tBZhBh8x
dB+wkqWxlVPopVk31C2Nx8oiyYh240DUmmhfHgiu45mwF6EOJUTmMW4aoOLvVmSn76KpdpGojFe8
+mAiVxcS25qYteqxDme1o4IWoKL3NVG//wGZTSXtWRR21JFx8WZvKOPWOtUvYCl9Z/lELUcmty59
GBHJD+qhe0x84vbOS7emUabu+QBPlspQBO1KW5GXHddw44tLoQHXYJsiacBwTQmmfA9FXoR91EhF
0kxUmcev18X3iykPesr9lzrKdG0AgPEUK+mgqveKPjRg79nDGZ1xwakvqQLGFrd+/MiD4n10t0WR
bhUHNvWAQ9eK0vxpbyHmv3TbLuUn6Mv6LBzQik0ayyCkxjWdjGtKvixfMyGbwIoDnVlyL/U2hNtA
HfTwdr0DRBLtFwLnxcz1DGgEO8cMBg+crOcD934Vz5vA9pbtLVv2NOiRW4ppFU5oiK4bszYfxBBA
lJYJP9rdxlm4G5C4KUMKNYAbOz8FqmzznJnFIk7ge/cYeTech3qIuzb4gH5VvAqUZiyRIkByxBdz
BhWFj8laK3Sn5aT5T9G9D7um+EjtDp/zwAVfTEzsPYXp00jXLmzjQWdXVES6liGUl/KpCdHIh8Y1
JEA1qv4QkYt67T0GIgyVyQoN5acBEgcxX4OHpJh/prKOId/A63mgBh4+xnUYiZ7xiDMA8fTZgFWO
ArGt8n14DfDmJAB2Ryktp61drGq6PEg5z0M7V5xQR2DbE/r/nxEJhEsCpOndBIKSShJ/munDWPUP
JMldpxVAPmPHYwKb0SdrZgECZOXnVxcFg+WjvOzPqRS1HVsOmwauu+zS7yLIMZ7SEG3FIQoiXENQ
2mr3MHc4TwxShi9e/0ierrK8esXMQPgxKtKyxAEO5+Iw1A96IJSRFdkVLdMACRKMotSd+5PnR2Wa
T3v+wohyf5RJCJaOYMVWcTbDAkzmXzQsGa9nlQe+MT4qJ0yYf9mWlCWa3W0bP5UQvi5FyvEJNXnm
cy9RItf3z/uQ36/6AS9FaHfydMlPE8C0Y67VyZ0Eq8tHqEP4AQCkjMz73BV6sF4stZRSJyBwu6Fi
be05JFRfTv6/7LIq2X5ICzTg8N3MuyIIMajqWwbCFrRbM3FA1EXyik8XQb6MNC+PDaM2oi32HQQw
suCLjgtbhVuo4D0MRIFBkRMresZQHmvh9KWd5JQ21UTU0RFQnMouvQsG0IPZjLAunEyO2eqJqL7R
kg4xehKrOJNNmkmcAtbzjmf5Wh+/jAL7mGspIhU8EU1lwoFN1jyY+cysUdrGpaKr7AuONt6D7Z0K
8J1jLbGBKbv8GMaacik2aZbE1d5EDztu+sT9M+0ApaM5okKjYC+jynn40PHW0QY/FXZAY+wlDBVI
mFdcdfLcQ28iyRhDJTQwNI6rBVYpHPIrRSZAJUsgGm2ovMc0cPLjUGlrVl26NTebUgZCKq3uOp0l
B2koCEZAh1GS8GQBCTblHxckIb1SXuF+7nhcq1z9RO3r7lCNKgqCHszJ67CiaYGBGsH9u/xG1XFV
5NlG0SyaQy5BIYo6/h8tnpGomUGe3dTMuxJeX6XkiOpmYx4UuNi1Q8Vvst2x1sDOikRr6I9ZnLr5
YCy72A4Dr3NURrurLTCEkbQJAvP5/yZ6zE0XQXrpSc5Lp6FSMxKJHuYWtWnAdDjq9gqYzeldKYZL
JfA2PQDJXshsFyCI/7Mnd2RMcu1v6PZBpuSaoM71YH/x+x+hkcdMUUxPd6T2ElvfsDDjdGss9qIk
8P0bS/TTi8D6VhePQc7af2YwFQLwuIPpfyHHUmg/g/5vzk2HdGimZadwgr9B7oJ/bMmKONrtbddl
BW6q8DeDCBx7dDEnevyZ9DiN017iHAqK8DoJegXpU/8my+ehutU8ePZRgQDSuAQd6cdrnCm27+7i
oxlnXDYktpbuNTvrLkjhWAGmv5ZRIKCZC3gDrjVcPeNF+vGCzLnk3RKi2p5rzl1Oy093TzWjIQYa
tJl9MU8dHg73awMWpJyEQcRlRw6Z0T5KFlxx9ur0qjTSsUg32059qHXCjGqddC/USKJrj84ZdnEi
FxYhGuRXFUpSVxxtIFojzJY2d1KIB9crYCcsocFKlBfovuxitiufkPE7gCYSnmzHyTDYBZbP34Bj
czmcXZVt406sYYNMCYGUkRHL1J0pG2sr4YBRDPbTuWy8tBMXocn6bmqV22NY9E5TIqUaTyNCIYnO
Vnc87cJs5hs3CrH6/mjFcv+tT460D9bxvWcu1fjO1jeFAr+Y/p8d5ZYJjcRZiPmWBFOczYOgi88f
w3M8XlarNGvwtGVOmSOQlLvv0rQJrrMpAkdUUQ+1R6mBuDdTGhZqu22YwVpvROtvDmNo+EZAM/oO
iah1IcMTvLZ1Wbez7yZ7qHCwbnwmi1b0mlb0T05JQS53RRCydsGrT4EO1/OTGCiQjA3w2VnhU2K7
C9m/DtJiYcdOFkdNJmLb/bIdWgrs4Ho3ccRQNie6K4xVoMGGw5wSpQwLezxuoCjKyRiduymrAEIG
lnTwSwcwvjaWRsMxgSCtZApP/H6FOqQtTJjfPgdFavsXHEo+H9hS039jFFo54g6LPsELbcO8iy1A
ZDQnhETnUCvxpKAoN128O1IXpCUT6oO0ceZPVN/+zyRRM380zo149RhYWtKdjJXWwS4kstSoev+N
IlFBrS8ILbYGWrK5bQeAgm/GtA7iNWVc/m3bRBn4Nq+L8HLA+9ESyViSdrLgXGMZXTNxoexjAg3Z
EuIk7ff5LM3BcJzHaLwFGP5ruC95mIKKiK4i1A0YSvd6K0YVNFIhq4p2nubt6FY03cvEbEj1WX8O
ObCGJaXDoUFCNYMncRSUyBRlNDsn6fMeEMv5JMjbLStyg7wNt97tyCJ2TovNWz7L0E9FcTMiJEOl
v+I7OKkTGpzu2002nPI/mfK7Fpe1Z3erjokhOU+jdkKwbauzi3gr7pJzCoQLdS81laPLb7fGJUhr
7Hl1ZxFsRVpa1E5tkHsMcusVG3T5ikWlMp0m51tQ1UoVrZQ76W4jLeR3EZV/n9l5Cq/p7DL7MAhX
QzM+ZjQrHIrhoZKb4URys+xeoNsf81PwD7Vb5HEviyuJMmTyJH4nl3Vm4l+cQ3XocGF4qVRFzF71
lHd79HcJqPds4lsgasuo+DT7u7pYvrgYyu+raVzzHnzGe+Wa6FEGF6erew20YPMvFkhvb883s3D6
lq/hwFgMBGI/Yd9JNNPQ60AzHJDzMWGUUdwsneoK0HRIIdedSrWyMqOc8yro1nQB4/a+trkG9gxi
TD1J/qQvPHdKaow1zzYXg6aQuDKs4GJh6txTzOsns8M8OEQBRLX1geeQSB3imCRtFWKZo/DDpdrv
aq5GqCrlXM097DoIgUqISG1W6gD0JZIpxWf3v8VZ7tJu9i9ZcAUfquS/6Lh/7j6om4Qp0IGic2ya
+47VqnxOlxmQkF6Y94N+c3SCRQbSH1+z3VDSXvnVyXu7jU46sXMSP8S8LrGp+rhSwbyIa2Pj1JBT
enI736i5xXLD9QkAypZasODqVnu82Oxyys4e3+0omAqskvcGRMj5yzLlIniohHXuE/x7uj1+qiT3
VsGq/DAVg5mKK7q3caZCtrP28dk+qgBgqMlfQmborIAGmxumZI0I5E29Kzjv7DLNoBmkdCIDyBYQ
KzfzrGWVzDpsjx5j2WVl0jp2EUlJ9nFM6dw8MOlE3yW1/3jo65ARyaUD3ygSq0RdevP2aLz9LlHU
KNRca4UmjSOSQ0lVs/z5o7GRCxnjPCT62ZN4Z/z8P2FWt+kCMIdM4IUznUMEk0QdJ5NlG9c4cl8x
/KFPz36+KyVsYW2bX1nI//0i5IWKFt9ga2GFwEbJTe7E5/gbE/AGiFiuGs2SXWfhYmAxqDvJ3zfh
G+izXik1bgP0NlCDo7k2jIKP7rV5LdPE2Rg2BRogGYSu/Nrz3wYeRMNqpfpW291H0f4PZajTKuW3
iNSv+enItCPtLNsyAbsw7IamfdyuzjJKg02oNiAfya1sNTX7lClJ4ttk8W1OzLO8nbmRzzON1hqR
1287VaG9lHr+Jb0iS0bxzdT4OAlDM8YYnmGBtSOYKZU+sMcl8N2ov6GdXh5TeuDyDGF8TZrdLT39
O/z957VXQ/SofhrXObYJqIX+QVLmmdilycigKT8DzVhBaY1T6lsrL9+/XORPrqEZMa22t94AOwKv
EacHZAd5x7APdT1UuHSpX4OP0cnL2IWMIkFxFoE2wg2QY8pGIkRaxVarHzZXMI0S7Cc709pMViBZ
6FnQZdKzs8OOd5HdBBVndJbe3yUUqEVMkQ+1HssIm43YQ6+6aTMeV0RDo4RVjcACwhqqYCri7WWu
sQknbWnr9b21xrj8MyFsjrPed9j+U89xsFcQhfj1uFdeaBulEiuzmLwSX/eL+aWgebaP5J3h0NG2
bHLQoHF1pGfNl2+mDwjm2UVnZm1/Z1scXrFdU4QZPRW7RYT8XUK3ycBMz1PEvjQEzG0/xm7akEfS
FUnDD7WpN8q0ML9bwju5FZWrYEgGAXw4XzXyOC13cXozZi8tqaDIl3XbF8E/1ZWbcaRwbTj+PfCi
H3ibJAN1zTVMMrg1XTDI5USvxQ5s0SR1K5nPDXTdcQmSdL/tABjgQTunqI0u3RSrBJMj2uBcgpWR
tE3OGXFCdPVcuZCXQDRB5ZL/Q/aReAqB5qutm2YoVXVAM8SFRfgvidIGgMaK0mkzWxOsicgsj+M8
YJFUmQvjT86sL7/xhUxLErp2iL6aI74g4CxbgyWECpOZVRQ4PIb9AacKLRO9AqMFjJ4fw3rco3hZ
139LXI7uXePkyGaRaogygS72FsSNVpRh1UjEOK/i5pM8PUvfXmqMqAZxfvXq//EdXFDPiQ0cd3QL
gXxdhEf32f2dy2KJOsisHy7eNtTLKmZ7gmfnRaGIy1frNBqPAaK0YgmU+/tGCkj5RYf3Zj95ZqaG
K86e2buRAREAYseEHVxxosxZ4W7pNo6nl1r6ptd6Fa/IOfq2AHiwkXKgeOXUjOzWlUae/PhYYU+b
UPXz7dogpSITtufVG+pSHwTgISKmlfN/ldFStKxaqDTgu+rQn8UYbqSv/ko2B8Ik8g1aZjuWuZcT
Vtm1gfWSK/R3IbU3vqPJHJtBIuq/jRJPrBiwxQGMJ+zF21lI4CBMXngZkyxFY2KsUepcgMQT3V/e
2JJfC7xL7lgWtGJBhn9MOoPI88fhU4KcY9s1CubLY48aGhP0L5ZtC4TACYwL/0HPOL0LzwDR5XPu
6VqvmuR0Bt3QPEOzX12K078QVNdlzsPtcB5D2DTohkYEFw1cbZclmaMGGwikgJiwK/WvHUXYCcn2
YlCOTcq6JvYWYuhx5J8EOaVt/Yg9GF5m2AMUccCZ07sSze8cc+Jjgt+kyg7O4hysZAWJ3wx/etj8
iHwz4gP3iVbEC1IjcDMppmjqBOmjoSwXZk0S+wKSE9LVzzU3y1ral8YTY0heweCzLnDleStm7fN+
nFAnSE0hBAGxFnXsEmJ4FVP+LxQNLH/HVPrjtgMW3Qc1PMtGYXrBAIOBG04luq4lsTMNLE6zgrRp
3YdrTuSz3NxzhELTj9Sqm4vS0NkmkE2DqbM+BpvCN92e1ywDA+AcyyfKpHSd2kr1yHT2At5pz6g9
+4Gt6vRtMAy/HeaTcEt+KNWjICCqSVfHQrwErYt6iUd8wmwTvxftZBoQODFf8xnV2HKj33Pnx12k
mn/82VOF2d08yyBMy8gv/o+UegyyWj9Lwo/R0nxI7DXIyM5AEbm2bKOZUfE1Yo2FSLM8xqA/yWvN
ZKbiiJz1xXB6YTINrIGvZ5lX+PCYfaaQaOU+mGsTnOsKAU/9VxZFBuhmh2MoQpheCYPgdNLxC3Q/
V7h50YLx0wzSJPqum2VZgEIUK0ld9zZqk5YHoKRHTreGZYEOlMyPk66uzskIKi1Qa26WU3hTxdxK
emAK4SKFlCkq0WCIUOMrvoNoqKrAhNPNmb1N49vuQhq95Rq+WZRGhZzApZH2JKloW11V6RKmDG/R
47HDgv+T6mE/SDqVt4w5ERr+ymASilQY/zpBMImk5N24SRjTe0fYyC+J4On3q3a++R7Jq8shTjIt
uKrk392J9dpnMLBqPqPfQnk4pZDswHu0XXBlyDcPeJkf2qhm6VUtxoD9o7vfllXUFMolHVL9Rheb
iNRHcvef50Sc6V2K/X2WrXvzreX7Hr7ZHscSYS5Ctozdbiw3JowyuBEjiZm6xjQhhg5qC90MGssW
sDkxL3rf+u28phc77ie+HAo0W9AujiCH0Sj3UEVramm7NYx9YSHpoN7NT6IVvXNxwlB4DqOmBvBg
G0ZykAk77/B3X4RKbh8hq26uyVpMdvL35/YWhH9Uox6ABjRWhh8eoGsTrxseriAriROF+rAhhGMp
TNhmv8NPHp76bNHURt3ZFnqYTnA50Ktg/CuDTrsBazTmzCJtR0JO6XVP7q4kIdW3BQpj3m0zJZrv
SPyNizCYs7myBSMHei580xqo/P3RDsn9UU2cg5cA/0/o90FcNpMZ4+50jfnYEv+HlaVbPbEKDwxL
u/H5CKSEDzkGX3XDRRf2ppdYhNziZe56QG15721F8VHUj+kqezfxynFH0LfrdvCFhmLgV1B/eGbZ
9emRLXlLWH4IYx2SdWOWYqptNb7PZZfkqtFVFzaXJQM/ABhVTs3q29pkcDgETpZ9crVt+72IAO5v
HGp15n7QwfxSGGT1Zuc88EC2YvsDFVqEd/SRevrXpG1Ixmv5AnvnDa3DBLA+OuK1TR5Jo0cR6RR7
yYMCntkBO24QRXP06FhxampQ38p1xPfSkxlgk2j3VzXqca8Q9FfwewsJMzxdExP4va011TVjyHA3
6jmOLI+BsMzcyW9uRl1RgxO+vHL+cQAumu6xnhIZe9+LAmfAPpeMxRgkrZwVU8CLozzwfIO2aLq/
ddkfp/Wmhuzy9f4iUPXLrqpBK0vnATSgeD77eZVxQUq79CGdwEi8EtnIxAEFXgOLguVZUqOGooI0
Brw7iXXoNOWDFQxfJf8lT75NByoqU2BKOzrQaJeRzBDd04+YzA6KjtK2yyJ2P9riaAwfAXNft/OA
42mjwfaHKBqXp/ucySCGA7kM8HoIRMaAkYcg34fzraoSy0rK+ZXwNziSM+Gm29BtRbse1fQFMWS3
Q4zfXi5zy+i5SjJlJl35vFUzj7bUO9mLRDpAhAgHkMwp7HSuJ8YZFRgQ4aiAXi/jXLkqHJdUBQWo
ex7tPd57+Chr+OPWHMFcpcJkvTEmbRjXM9cGLxzDAaxvMd0cFK1mRr0hj2PP7I+2XRMyq0nBDQ6w
9oqulOz7JnPNA3bAAcjq4gusRFX01XWZoD9VWEq2XdaLAcGCI2SvI4qUD4RTuYyLl9cTHZHd3QZw
bNpZFwIO17h46v/iFObg3TL88Ueipq93O3TlcueGWWTeame3j7jlvRmGJ/LppVMrR2F8SDyiehYh
0ozh2o8MBptU/HtyAY+i7WWH4H+RByslk83z6Dx6+57UxwGAN1Tf/MStPCZy18rfjRQxceFdfWaZ
pyZZaoP77y3aDr2IxGb9DP6BuO5sGBIIXEV2sXLd65n/pm3PMtXkQvN6L8XcVt2Wh7rpyMQxo42U
KXEfadGcS7r0LCT+uShrickOgkad/mKAXvzxkbIaKRYimjIvs9rj1FiPqOflA1hMMFg0wmAFABt9
XIK+O1wgGGSHwhdpRwLmUluekjHVGiecEc/owFr+pKfEzz02Hr7sDe4C9hywmmH2mhWmqg34Yfnq
m3s0xP5FA/GtvEq0t+iLVfodR1JwFcihUnCq9CjLtJIUBXYoIDNa+5rGRtw0GgK7uQlNmX/3kiNR
CMhmsj1w+8LEixuD6QxPfJXgvsWJSXZ7ElAWmJllSPCuAdO9tMOJvUFuvz5VM+9recZZd5f6SIcL
S2mKZbIeMXYBX9jM/vrcOl2+2KUdZIGh+yQ4/l3mMUxHu+a3gzJGLplUy+QBrEmwRLFvC14dyVhl
X5DHf0xJ2zXhaCA7wUELYbj6ig7UUBrhme75dy4wQ3Tqb5KyR/Yx5WTn1HzzMHMKsIyS7/dihK9k
QUXITEz5NQpsqaEFMnjb+zFQVt6KGXgAAVenCX7M8UEhP3gCtLFuDx5W3MKqqhdkyqYD6ZU2Kwjb
h6pIPygdZ7Fbr/VSWX/OiyH3nQN0SWesA32gfJET/55S0oACWeB6ln0Rvr30crbxocEvzR9MO3Hb
DHPNwHM+daCH6CW4rzlOJTxYl26RWQis46oIP2p3iqUDFYCo52Dd03pIQdAqbQBcmpvgTHA+SYtP
7o3p6DFaTfg8ItpysTtVDM8WBO2CCJrebBpY+A+NxTQ+sWWppJe4p+O1fL6FyYN3gtP2itrfXsKB
u9zeuOjYor0f70apqxyMwu/fy9iiJNMl4NJCrDQw3OjgVwwKjO9IawhMbkXLgpSf6oPV56V7nAvq
/ukWBqt+zb07zQP4WwnBOkxoBNvY67oAqrFJCVgFMLsosQarjrx739bFlfUvdaD25YhkX5QDdejm
dt7872T4ZE4ceo+6R+Prp0+Xe3koejMPNrZWelUdmrfJ8yqe8LgWdcj5uKoHacd6rkvXnPZnYjLK
Sd2i/JQq0eGaalq91hjeXDmdT0E/lfiepOWEdB3hTMYgNQHSqoJ5f0Ntt+kDONFvycyreUW+hTjK
+P/4ADWx1YjOM2cFtgj4nUWO92hd1p1Bd+HcDwZ+fieVFkqycpNwAQgfA4RKL4LHUWdxRSC7pCxt
9BYLic6E/4HFP0wURkHnTTWzmCMOtwHRnEwBClqVPnUIdfgKuLw+k8dhAIfbrDf0ARS+q6sjPBlV
H6Qs+v52g3t3mDvwBK1C7MQ5ye9E91eW5jL/44UW94wHYLXexXqpBnj+gD+hB4O+lhefLjGkWq+8
4LrntLXL+Zi6Hz4qAttIoG60/7CuWKUVLLhJFF64TJ47+gx8DDuFlNojNkA+oKYR3CLylLW6CbD2
zvjxE1kysOm2WzTF4Yqi56PDTY8xj2AwJW/vUHXibcZQ98h6Sr55RUDP5XMOeYZTaYN4m7K0uSIB
qLBMvx5vVB+L/0M2G2iojLiNgwJRU6zSTORhCPYvsrUu1FVSGN/g2z+csdnmT96fnJECmK2MdEhF
LmJgeEzXl60IpRzY2Ju7YWqimjjQ0YwK9tqcHrv6WsikrHOKnw7GfmHfL1TMhI1nIZ4zvLvfl32H
/go1LqdGqDkNb6/nSNRptLV49FWfaAQ2v4jDZgQErmcQmDWDvMox0ta8ZIvohK4kRYVkmQcSBmCY
n2YwPrCVSVKwlTpZu5oioQrdBYQOR0YzSj1bFN9GEOnaITHiQlK+s5IVcP9CGylvZjSN510ADzSw
dXUdQ+CiQMWz3jNJ7Qm+0PQ/dr6/cY5rcilRWibsJ4Rs8RaOLsA6EfhmC76P539Ddo6ghRgemS60
KNDquqWHeXJv19a8C4rgDAtPXT+bBKsCa20pvb9ZSSbmTYV937qZW8e8kHWvYXkb+rKVy1FJIvhM
lb2IuMusknjNBEb3Eaxa44JHa1WOFkqYh/1gS7znCi7GgRXB4a/RS92kVCYI4J4e/7atsOOIf+Nb
tFRNsOsWWxiKM7xnuhJmjuI087pd7If+Vp39m2K4Ci92M1t6L0zhKtECsTo+m7ASY5qy/+YhsW7g
/tPNbrRHnDZ2pFqze0yM91Ky7uy9LyVWLdGrvmMIYK8z18FcZZrkyfNKZhj/nROCcf8/xiNG4Q6f
lDDjnDry55FdkKQAhj/VrRn7c3J554WauNkpLRV5azzVFP40qG0dpRAP4IkFSNA2Ox6dEdLJQS7t
rYSmCaMuzqGC3DDJSTjV7M1MjcdWh6ynBM6GEUe4py/NSV1a7Tkb5h+o1WHAX0bRfaaDcDg7T6ne
h/8iWHOTLkUlklkD+YwGj6yPHuf+SnZouFyLGAiZeuHsyBnT10WhuM/OQqt9IntSmH+Wgvhwu8fP
kZh4+dfjgVdu2oMbnaDZo/oecnnw9jsC4fo5EKM7lmvNa4iLeqAkquovKTllg4xUPb/OSUtP8mmY
1rBgKlijZR/4SdpYhZgt28YFMoFmhcUJk4SsuUoIKQIA9oO69PY9J0juN9WXP6gqlWnwbku8SsN0
mNaMK8mHMVmB1kufPlTuf/Mff3QfRMAnXjtRQEI/13ntpA9ZRR6IJtOLjyftC8ishqtlZILdr2qJ
QZwNC9iXTS2bLGEt5Gqi9db795I9iVlOiFpOWdaO+2zjnnvGnWBsegcV7wGl7XsQeRGfBAlFj2x1
NxADWB3tcWkmzMwi9HfHkDte/glor4C/r4AxN3pnlBARzG0cGluE4nHWR1woR0NTHSmtStxJKMJH
1thgTRSKG8cZzFMz0ul0FQnHRX3cxA+i1mwJVOZAWO/yPU70ag60qbGi/gpdDxhHlGKDh0+/Y2su
P8LPyZRy8u8cn7rKMZcRQPFBF5olqFz8p9p2C2wIKDDt+of5x6fYiK8rznMkv3jOAFxXlRD/vr55
J1LKf4oSg2QUg8hMcO3pMKhQQ4MNAmjOEtYe0/Be1Zvr3hGrsn4V86+3m4XzphfScKbGPy+ttIoT
pvnfpP1hDZ0lL57b4UrHA+PDpH1eU1DnXxAbagnxeJciSMCcRiKU97z7V9Wjiua6pP0ASt9L+tVC
X/HVZAr/SgQtRV/wfojvtH8E3TVMRkbU0ZUSWWHbjY34EJxisp94v0bTggVnfB8Tz1vg2Vd6Sx54
VUPwExdsf7cSsAgflDs7h7RSwqSXyItxyMXhjS64MtdSG/DM4PlbuZVw0uLjoAwHvBN6f8AZHLki
HLMEw65Nmm4tTdJJpcPHPEoGuA2CLy3DQ2meuF5xkOM81DQ2WfOOXbXDgYJuASyEmxcjpnRxuvQi
1ISf0bVL0GevLK46mhlHBP5A0w7hbdIhp42hibilFsEU42Cy5uyfW7ymINaDI+F7xeF3ulyfSI0o
S9XN6bT1xiHSZ68/45tZaPZlUk9Wqu7m4CckarEEYSgLGoTU4W5uAcWUvE/XQYUTTwQkArX6tlMD
TMn5cOm468/qSUc5Bshu7F6wXiCTkLAbBBj7Xqg1UpAFYU1idBlZ3RARBkJWtTuF0/FfP3yNOv3Q
fscokBe7S7YRfMcPktXazRwsFodke8/TkiTYmoqjeCYhBByxf/qtJdNT3l265V9CU9yqg2waNC4f
530imO/HlgfFoRHIJ7KM1Npbti5nplDDofnZ04SOk180a7yyHiNfEnr4Q/G6/ma2Zg38Hs2/AeJ/
DmEmyXwjsfHCxk2NQzrOtbP8sMBxnMu1Jqfd0pBTbV1n2y7wJEjZ6sEWgb6vRAJdXftL07+SK9g6
Iq2CycKpHTLdr2lI9QSLfzi9RXwbzfHL3urJgmzRfJqMeK9WCcJu1lGWMlHFHtf/OI/L1rfSOzGx
3lwwN+5G8CAnsrfDTfeoKlJzcminjSxTHYLl1jdRL9UuvEGfHPUGVJU6H32Sdp+IBi4xcPatOjLn
ai6F0jibAJhgKRZac1wdi52rYb5B0kTkYP0VvK+lMqu2jXSXwuI9QLA6rxOwHkiSMPBmRFJfzAU3
8X+SeP0D3/RVLij4kZm5ZswfJikKu2kOA+6DH/ewhEMiO381nBrmGHYpviSf5Ao+38BsK7wHSK25
naQ6V4qKBIcJHzYe4jQoRl4YFi/ArURRrpV9cGPaa4dDk22rJ8ygdZjkZig/LeFfjw+X/BWWzdTI
0h525rZc5uy88uS2o77tymW3f9ONpVvOl1uLEJrfGI/PGdXR8ZFmrqoPGuY/cpK1dK4deK2HsSDF
y5UhExrPPJaB46K4TE5Rnn0ECtBmQzzPTimJOXiLyeJivTAz5W9TOl3u2bI1heB0uABJas4bVs08
I8mkZ7ffWedhdzC8ysCc9tu3JUQWWME0haW3Qr1AlmWU6KPaSKQFJg5oCJrcdbSwR9MMOCjgboA8
y1JP2iC9YjGi5+L8wmGlIY7i0L+WXRnlYABJgn9SPIhIYhB7GI19VKsM10x+3DOSIbgekNa0goCI
3Shaf9dzxkqtkN0Ovd/bzgLbcsDDm1AkF80EYQM8np2biCFa9XRDY/V9exUDHdu4cGRSemlAfX/S
+6uykJLTodRg9FHlCGcIZSjQvQZT5ejS4Db8c+/+uSC/j7mlugSNeAqGIQSMxNAmZsnTYuFb33bQ
KlBs3PEGfvehP7tpZ/lTZUovyoX1m+ncF2s/kkL0FTy2jdZ+xx3yLRKnUMHTban2aFr6sJSK2ino
JrD6UvKeDD3h3awrclU1Y56L/2X2NY3klvOZQF2ChFDJdADi5XQU1RNto10vxykginOp5GhDFS0q
NjkHxSrR5DiXJQfeMcuQcp9a7TMFX3qi510Ev/oTvf9og9npJW8oZVYJGE/ZWWvafYmCGzMDuNsp
WTJqEncd5QR018sernWcmmSS9AbFnCUF/s1tIrF9+A7OXA22MzP2XaPsgu4Yecw5kEnKt4RilZJ1
opxrp9s/uQLuXudqMvxE5g4NqyA/yk+sxa8V+tHVOQV1j8pAyF46G3zy+Jd2pCcu1nHQVJ88SCCY
847DE6+/AI2sMBrRL2ohNn9HO7mcD2qVTV/8Un9nM4/+f9Bj8lP/MB6nODnSAys+a9ru9uPXzTIW
6qM3Bz1DZBTClaQ4esIBhIh6z3c3FzQYcZljXdLxt0aYykEDGn14w7I3qWVipNtHP+j1v6qDj6dl
459rn8KtncfVSBFcTf4YNg2uRxZjpK6M8WkMBVDKleDCHlJg3S180JSzHI/hFuHUCuiWAaGOxv9S
5RJEUZWrUGeuyWlJoZBP2Kxy2/n3p7P3GSSXoCwcd0gRtTNBCqtcyO9TmNBEcEMlKzlmJ6CEyndR
twcRqXoE+KXZq+HgP9sCF4oPESZ9tiAsVJI1Zi7Lq3dyaZgYksjUpkcrRPTe2javy629E/y62qOJ
Pd7R5V771XIZpwenGsvzy6Jlh88IJLxei5ZMaMOpv2sdBqXLTN75VR4HdWvfjlW6UY1jkSkGRest
6nX7WNtVmWrvWdsi9/ya49rh2mM4j/UQDxCJhxeiUlKZyqI8ISCvDYj2JT6NNSp7Al8y11sAtXzE
W7QkjwTr1V6e9Z6H2gwyAMNozcJRjtAyhrTjwdZ8A9K6QSfXxWN8ljH/xToJhGyE7V+g7Fs4UAp4
zANeQW9l5kLtNhxtg5JIOlOvvNg6u+E9zv2264/I0Od+eS1qNUuBE3oAeSOBuqYP6gSPXKgqPZRN
r/479z2NwnA4Xje4rwOhr7QK4kQM4+AYLtH/5DAlUGgn3o6679/TDVklR091rU5y5HaaXPrKOFze
gXViOMPjCoSFZxqT55zCwS+1dc7Lsh+4pmCNg4t1DkflL0ceUbHHsfeZuWleQMm2iItSZc282U4V
xWlAzoMB5YFw4mbCBgfzBK7U4H8AdX2cpiU0kyj1kdxG6CnNbm4Q5kQG46rMB/hoU151MMCjDL9G
H2jCnlMX97scIVtaN7TGyLWWG8hxK3St75w2uWlm9bf0BHtRvyU4/oCiZ0smc3fnlp9M34VQgIBC
QflG9O4/d4xN/weF/AF8D/k4jX7f2C4eqctSbN4txHdvb5k1txNcxIHAe5m8KyTksbCIXH1kZgni
W8kGH7/qV/waDM1ontNheT6b45YLq9so/yr8kD9W4LeQZBJ41URiCxTEezAJ8UQ2ZCP3crwUrtSU
jca0le45fDA9itHMKj+/9kulb8yhAL5+z05xvIGWB1P7OBX94Lj9KsWtTSVwyDLLF8w0KVWTlH9k
BopF/mjDlTQzXwVGalDbF29BfTj1eMZFAZNtickEwJvF2Gy1K1WItTGTVc58DdTNBanNykwix3u+
IGH4h+e7WNQvK3d3up3yDSWckQn0QDK86gEO+8u8G6ke1UsK/zNN7goBhdTFfgQUg/yFZNh51OSb
mMQdK0NZbn0Me6B+olx4pJuth6cH1B5yA/a7GVN7dGvOB/GF4J7Lsw3Lh7wlGMiHVphFKwWG+xCE
18Zp0MeyX0CQJE9qDsoTMzd9EELBAkIvihPdYl2jOjPmTyUVnW1oNF+cv4W3cnEYC3TJewM+UM4q
ZoeHJbROtsliW7JEqS0QL02vwinNKyZCNDsXdFHlO2tJia4nZU1BzX46MfhihChkQV/DP8FeLWxC
unA45YAmqaP5chSYQNqqCexU9yF6GDNHoID2DCzNXQKQDpZcGVKs0RB/NPyDBh/i/1+OCyQFtSzl
fooU6BtTF0UpXgZ3U4GjB3wgmGB0xXxVCFvuoVy1LqanJR+G+h3uVQlzQPwElqhys36MjwN4LIgS
xuUuzvlGXqR1WUkZt+zp0B3Oi9HSm79J1JscwI+g5fc7khasVAlT83cVkv15oV4jtQAufmiKL3G2
U45R5JbX9wBc7+s8Ao1nBSV30C5m83/2z6Zbm9bQyL2uBI8q0CiRXITrsiSw7QOu6ThpVvKWRweP
wvXD6/6eThwzOzlDlVECcbcvFvS+iqxdAT1AzReI/ZFaBry5hbK/uVEhsZigIskm3fCxXfBG0qRF
0qdmKWJifOcCWMiOiTpBCyL/A9B0q1JAqPLVFaQnYfIZEg9bAacz1/sBYCYfcOCYx787HutwP79X
y335+343euQqFkeiesCk3ghriAAJNIYJv6SF9sQ0rreC4JlvXi1F5WMqBuEh42xYP2E5JkK6L/8r
SgMmnfuwxPeXDJgYY7URcGB2gAtblX7L9lXnc+unb/XuVVi3YbAJyF3b5olMkwLBQgDkeSJKU7P3
AJBPXPDcMcpDrYIcNYKxuQ/qmJAPFv9mDrtGdRixnzae+YCT8lrL/y90QpspHdihPnYkzQN9RGgs
q/eYp+iYjlZsfgaYH4YPoAtWyTtj89E76/7yz4xrm6vsDaTDIpqcBPkNCOE5jchegiwdnzqheTcZ
6FedecKPQJjGUhM9acy6Xns2sJbJmpC0czSg94Mbey0Gjjry48hk0eaD2PcGKaUbvBQhHchNoLZ8
EvAc9NyTK5ZzUuetW0m+SRhQYyXn578uXhkpqexvuxK9J/5H4Ca4eHs8BraIvKCqXQyTi+j+stE2
UyYhnBM9xbGg+2N9DbpL6mnYNg+4Qe+FLkgVf9j7GZ25IWXGh32QlDMs5SENurrbmEwNVQVaNbQL
020I2yeF2OqAnSQQi9VHQrSEkdp2fQooHKT0jeNuz/nwHaZF6JuPe2FjtMxi1C400GrvfWj05456
opq6ah0pzUROH/jmqeb3Od6fSinF+0UiKXRn8aFDEHKaDs15x+u50lUc1H9tQPpHzKLXrkjhKhU6
JG94tb5f6ViLpaANu1yXFknGymUDr9ncOcG6zxd+XeOT9ek+kTbidLAM8h8poil9LJCbWjKbozT6
XSmNUHnsbcFcLCBevbKgrOBWWAEG4LsUzceX5JxlaGzbyDxSTSljuzDVDSIpotcY9ivnB1SR69xR
XMBQY3AHWInnB9Ius6dgUzu74rD8R3Acmp7yJuPXopyHeEDRSCOlfS/rop5gZGal/YZcL8MWf1q+
8+EasZYQkYIpv21UnSYcrryiZMkM3eVNUcV2iS8KxCwqYiq8byg8PWzBOcAkfTOu9Wt9jaVSfJjw
xjaIuHOuGGanTYd7Zln5N/XTW/qN5lshcH33OBlQAzXGTP8rSH6svbXO3//X2O7s4GmVrsR52SYC
SgYvzqdSKPvzu0EsBHh06ATziifYOG6daQyqY3DGFkRI4nIJaF7bvQAb6t1hQGhUHMyrtgdQuknS
SIifd58eOuNH31yZ434pwko57BcltiDQlBpEurriyDTm3zc2Lf1/zqpejuLVpeRFlohjCPLnZp1r
SvTukI0hM6szXcL+S3DqPEGsYkTAvZZGZ8JIWe1ukw2WUpTL3DxygrWvH0jjcad8Rb9ACx/MsJWW
zJ7dw2TqvvlrXwUMsUbFo+koleOsRGCsdYeIeFM3dinpdDB1mkO13ZYExzX5UUPfSfxt0NwpaSN9
pGH7vxT4jFEqmwZPufw43Mhic0G1HxJzoLc0nyfoaYecaH0QmJXsjoXDw7c0LOB61gxN+7YzYZDT
YEAFgr8JBatz6N5O+yaPIiN1+ZT5uPwPTmMsbwxYtTjh/vLCGMMz0JzxHRIBIZT7c5Lsj0Bcmt4o
i2l+PRFtK9H2IH+90mLBl6tdVJXkOMj+AtK9tiIm5orKudKsSDdIbKUbu0zgFtUbUKxaQLntey1N
ghgf6UBA0DXZuVafCefSdWZR0+xnadEovsnPnR2iy7RQEwnqoVmhGq2yn2gcySRFmDHKggydj/4c
MkHqb2CZF1YIwfv0X3EB8RogfQ1GyAZMPk8BJ+NYVuSq+4H7ngB5a1pk3dgDP8i/I8CMBRa1d8GP
3J11kR3PuksCtlBkg7qa0kEleN5+iXlj/ZxitEF8hcqMxQhGJPseIwzDspEkRs18kHRXdmDltKZZ
PL5b70qWxza0Py+jQuaO0+128v6HXdBcGRlbMQGz0P59aN7sBhR9PdNYZGNaQF1zYFmg11oH8rQp
vFl1iiRno/lsNUAkAbuTw+2Gopdyj8Q0xdFnvIBWos3/zCLKQvYiC5mh2Nilp8fXfyuNOKuTQyEH
7JtWdz5Kw/yYpOxYoswIuWfr8aKIczsiy881VOEPUbISdIMR+fWmBU0GxUp/ic4Gx9r7CSTPua+f
EQ2xK2ICQjyQ2/tBT3IDEX+2X2fRWyOCw4mz+EaQ6OJlcPDhWYJrr2dTRaFLnlh3rAVGdv3e6XD2
Ifwnlq8A00ptnbx+aO5652YM9iJxjP96oIqD+XghjK0C2959zre/FcSThfXeoefB3tlQ29cAkl41
3kp9ZeBe+cmRoHwMia73YsyZvlznJAt9bYkWLa1tb2JXnyXJIqsOZ/iUJb6T9ZtEWmY+ltBrqgRU
IrCZrPwpQD9xxboB8jFEP/E9MgtdhXaKEUyXUXTyHXAimBkD4JX9cFBvFm18jblY47YGOssvX1B5
mL1F0lg8mKvska0LY+useSr0zLDc1DIUxruJ9j1m+jjpXiAn00rISM3/O3JDjAnSjucD/2eRRX/F
kKrk/mulwoKwl8YXxamOAPo0jCjWrGc4MHDWKFNHwQ/CLK8LeXkqm5euWeABpXTnAxQ9mJGwbXUa
6jOS0balbAv/YgbsBtxrymHid3lxrznaEXte6rPU4w9bMJA4RwwIKem4DvF0R/bD9EJ80ZMM9plA
paJh+OwGtGoTB7GLkdItLxb3hsdzytlMaH2mopgO7rcSm3VB4TM/JwqA9xZ8qF4OTW1YVodYEMcI
pDYFqTz3bIRjNwCrLzmDVMo8fx+0F5zXyEkWmNSQXeQL+t2R2iKoEey8Oj0Vs+rRLwaIbs+dAx2W
qOhT00VStcAWoq1FVcH2GRdmkSa8reENMfLoi3uj1jghBsO/0yPIVzHqDQcsA5ExfmWf1bOuFq/h
8wlA4igKLtLBUytPRl9FlQbLIfBYX0SeJ1P4F49Hp/mFkI6evIQ6mKCyKTWoX1Nfy2HwFGjMRq8v
AOZ3Vm6GtP6Ts/+mqEEaE3PO48dkcYe1LldUQq7VDTorvxpk2F65cUQZvZjuCZ+5GqpGem35Jq1r
jBUiVQLMVk5Mh62ZHVCTT8gb3V9agi9uUSpBcLK2Y1j/Tt96Q0dnGNYpLJgcoFtPL/hFjHQOliyD
hoDbknRSRBAJjwB9Q1YGsLxfwl7DJhL8ObSDqP83ddjPgxOrR7rVVm17ydZ3RLvNEbDMJDv9idlf
9Q3hcLDJ1jwFKv0vott9rpRRwK3OIf5q7ceEpG7rRaDV7eiFgqzPosw3TKCfRrr5mIV744FKqkXN
4YB3RWLlUeX0YXi3v6llpmTOFMTSvodddyTS32v+8WX5mehBknh/h7PMJRbbF5342CrbPBPFmxmp
ZVEivV/Fm3aXXpu2/G1E/rWDWkpsOi+s93sSIfH6SfvP1u7rFBYBYwGrr2s+iPiAND6us9KQUoRH
v6g46CkmaD0O3foECDvKVtRioV4lVscwtqkMmfJi7DE8xtoWDQLDAk52I3ZiKWFTuXbooEBkKCvc
fB4YN6kOZBwEBQDSPBmmQb6FZv+FfLptE9siq3UHQr71FKfb7JJjT0mZrGufB4enivIbik1sI+WZ
V9ItQXrSMY9KN41/Z4Vv+9UZsUxENZMXQFewdbMep6yM2lkUvWJM7j5TffoQjgiR6phmDtWTdIcE
Broz5upQf8cCbCZRF703CR30xSXt3EbWGeRlP5rmuu/HEj1O2F5KCOklmHh3hWg2A/8UeuDj8gLZ
mwaybwtIf4OWz522ShycKHI/KoOW6LRmS8NuorEL2sAOneVT1+HoT4xsMhl5jlg0ZIUWyomPHHon
wMHkBoEOrJSLZ6iHNAoOs1Oz0AVoU70V7CrrYDoUsXp48If/FVKuOEzOA/acVIiXlRentz7ZN8UH
c7Yohsb6wcmzQ1wycO6BivMZ19QY+g9z8r3zJI3pdgaNWAR3vWm/tOq75L/ZPA4sVEqTFkrECsO2
xauz0yjhceqmzFb9rzKJbGKUxdfkbsecywRg6TWKaZR6mk8XHuGiApX3aRFWe9w01hJRpsWPk7OB
A2i2nwcA7PdXkZnBy7+sJuZ6Dg/hxtbUb4RVrqD4e6Jw31SvvIOMSbyIvXe/lDnPek0gAV4eEnIk
jORoc93q9KDytkePdPw77CHnZP8bc8ncM0udiBz2GESAofXCIFdO19j/Gd5aZ+mYLUD3CASSTu90
8n4BPIIKzvBhAkrwXlUoYEXSMmRW63bVqjFnmlLZqtWWlqobuzZM0BHi2Hmx09OlyNXNYxMKoGOa
kL0myVFf+y6zTgVrCCju0e/HOT6JG13t/PYjji6gC07H6C6SL30J0AztozrNbt/myArSHcUV7rgk
6aGpqLoRl5BKoRwrPGv6+tO1k92NJ10O5GmfTVXuOd965jmpGy3FfS/tLaz4FLxn/M/vxZTEN8zk
4EeabFlN9tB3sMGKOlKQtwxDVU+xts+rS4jy79T9UIXbKVZ/NH7x+1Y3cHtDr72l2iOQmZSEfQOI
7wTG94CpnPNDEjam2H1Jr2tWoTfipUobjOUVW6Tn3reFGdnEbRikSxXkDjRo7IZybp9eebqTVDHA
YJEXfhABpTrvLVTWIS5xenhYgeofxFalIOaR0mBayf+Xo1qbEtflIK2oJy503kwObvF1lQOvNmE9
Itkf7Yq28lbMU2ClwWhVCSUnO8c1ABDxdyMfvcAvitDHZIQ+vmnIjQF2ZakRb9Klp1UVb9aPIipi
Ky0YBqts8GWei2ByH2J89ucY/Vr2Cdl9lvipoaR+aVSu4ZtU3xE2tAJAHff0IzIVjovay+L+ak/5
vCxpJNvhSe6UAoE6O8sbQ0i8zrZdXMS6wRTFLxqET8qdkrwkwJEx3pMq4FV8KwXIYX/iRTWIZvc/
azSKgbYuETxVubEtK5PPRgf05H5KDQY1S/n9qltfqUzZ4YR/jRh7hmGN6ca4j62TtcfXKi3cDy7I
ymTURTurQwhrSTJmo7GHDckNNA67NFQ8L2qcFT+03GX6Um26t2AraMrZ3sNgyzAhF5zCvZUrF+cw
ENBDlNwkyJMW7dwX+7njv14DEW3eWwWci1ObEDjE4H/U5smawD+rBy5i68nab9v6UpbVXVi8EMZ2
iyYc9X5ypVeWxjrHKY1Pz/tt6rCn09CIyk6nMTdjYw24lzqDdWKbwuzr5Azqqibo0ujpgr3Fqq5g
Bcuu0MdY0VeHZkOdWzq07p08pYAL8f5FRXax11r3nRxLAw+17y+WurpZQytjurxUSr4txVo+DCTe
mFaMdB444HOtiIIbA+Ghx1QMlxwpkFxnkXHuk6REtLBQGEtCKNZaK5DNNRqbMsX9KVN1Yzdsp2hl
Pemx9g26Pe4K14P7h+q7tklK2RkkGVYV2fxYd/FU4Wo4D2mxfoVzGTtWep2WsdQO3MpfzTda03fd
TCMBasm+85QGhtPPn7FH4hkGB3Rvv/f8GIgB637O9xF9fMu7zjX46R5QRuCGxNrIUfYgHkXz5MJd
YJM2KjDQliyccRjtfWBPdXByU839aJfMoB3L8IN4AOXEF/M3onxEkNRjjP5jHtUnzSrsqoqX3xMN
axTL5yGiXN14cRDBRRkhS5itJnPLq9IDCdf8gxB+S1qLrotp/cdjpmNeQC0cYYXTst6v0aRN2UBi
VcleSf5LCzrD/klAjkIDy+Nodz89/6gwDzEaaTtf72SlAmBrNkPOEILFzCcGy3EBAOZu++lteAGe
Yyr8edtXXB9/s/zIJuyt8a8GDR9t/X6Jg+PDEtiEhnWYwIw2yf0QoOa/P4t9XfTSmuLPUHD4VEij
PUKBfJ8eycrmkVnDEuUTtATazXd0vjxB+YtXZlCIOrWgyMENSChn9sa6FJ8z07mAHzvm+bSTQI3z
IcfiRlWJA0fKt+U737zuvjaZE9vhLEyAnGkaf+NLjKXWEFyDb/cEIzfQrJ0NHYUJ6QRaxDU5PnGz
ZoS+DwC69z/dLI7+82XBu2oXnjTzadIK/RujGAJ/EYiqt83GqHx7pJ+bUly/UZQDTRL+w0/hCVTF
YsoFzAu9qJzeRsqHSfcao+Mr48UTpMOsT720QwHBydWaUq1o0Rd7DXY6PUuIFjUVkv1qOrSnc34k
Ilq7ILsLyCVn8E46uQeP9DM+FSpgjhAmTP/KNyAXxnnAH0lZtNshdCjrlBY48S0Ds6OiaP5htxzX
kTYGQbfr2gjHL6LDVmDwIEK4dRHJoQgLXTFJ6bR3KoH+A5YxmsR1RSY0O6XW8H1lElrJa/GHC8HY
RWVuYS5vZYPhV8RxgEOb6LX37BFqFwt3AHUCLxOmMeWzDpKs5ENnlRnMLNOZ93a8zXrTGULgHtdv
WymBmqvoXqqko4nZOeamvlNqPbOQQg3OhPkCaT3l0TPM5dYo7OAGh16w32W7QLkyWiM85ooqYDB5
HzKx34qeQqIUAboMYN1jEtomqcnZDnqpWY5lJJ5GenCJ7SKTLVuqU1xJvTF+3mNjAIYG4+g2XM26
PLHp851PMVqrxIVHBOiGthSAWDA8XSfdOBihQhp0Xvo98LRH830Mh6dlDnzFiaTxiJs5mkitnqjV
dBJRM+CyrsXOMuXSkzmRKQCnkQyG56oEvPQROdffyT2aLpMNGSck3zt/8nZeWTeHQO28OVEBwfAi
CRSyYgw1SlITANrjZ0EwetbOKXHhv+IPo2ffRO/4DT88LIIesGVwKW3nfnMOBVavtOxiAdwAisp9
iNTJsI+p/nUNpGueUOro4I2toM8D8ny3pxuB3r+v6TSmBi0jInaQtA24pitwi5zRgTfWj2eSK4ic
WLJ4XYXjx7tsn1IkwxkBaliS02O26/vi4COxK2b7bA994LqUoFncaa73127knhwu7vqIk7HWRECH
UonG6LHK/GPO2wX1c+44WoAPQYab5noZR1o9aB0Lz8sjGZpx+3TssnN+7QhS8bvh8zvPr3CcDnGu
mls8xwA7NBrhGF5Fz27dxMsLWjcpVC7ySWMWZ+P7vbsiX53pQO9BLt/XQoe1okFrpi1ouzStKyWA
ptW8Avh68VUyoXgWHFE19OcAtdwilpOFXLds2App4OziuaI2ra9VBTQr8GbZmCxXtTLcNsoYN4wH
MK+IaMQxiiBOwYRP1VrI4bPSitYf2CMEJsOIYaLiZHU+RU9iPqhj87aJQrlu4PFGQFv2ghvNhLTh
FXxMOB5MPm+TVhn6cJdTrdsb6dTQ0imUPHoQzBQojm/iJgEv5TAJysOYjnUZvSh62Mt8HA9AG+VJ
zStlxl2ZRutbmQ4Fuyl95XcUOSIkdN4ZG1q21Vv2bdWo5olcVo1JvxOMrUXQ8PLIebFhtnP30HFT
7CmpLGdyU/fWszXMBMbSmdIumt8vkJX+1f2nh4XeMrl9YnoGgCA3EMzsIErJS+wZXz1mqN2zRXhO
ziVF5S2QE6vUoK4va3kDuXpmLI4CuHH3uTfxdHyFajO9v4SgCxJdzocQNRRzwcmJIiD7dujVay6h
sSOXJXG5CjEJIuLK8s+MyLbkgXbezsUcmJWyxfsYnE7OiP1Z3JkZTq80zba4ay7o6PtQiTh3/naJ
HNWJJmoUo+WsTZcd8Zuf1S0LkhmTxx+lnri0MuDnKNSm9VchwKsblSVX+leU1/VTvWpgnXERIaik
6jZCK6isEITARYRY11soP0KMtmWNKV74DJt/dreg5159P0s6jB1ywgtZO+qV7tHIR629bbZP+TT9
71X8Sap6nEL4kNS6L9piC3J4/22WiQUO6CjzDWP5BKZAsb317DEbs/FzFBLoPfaTVuRPI2NuNm4d
gBPk8s6RFazK9tg1A4fTZV54mVp1w+zhcmMy2QyB6q78Bw5L4npvPKsPYm6Dmz/gSckIiFTtX28K
MzrgRgria9hVff4zTEFeCPuioLjDKQcRLHKzYLLSKZIQJJQsoiLWMWHqigDcZpL3RYwmwuJiDIkB
G0Kkzf7ZNCAACr9+FGE/gG+JYwnpKIYO3YorzNILXC7ea1d9VahuL++8ly03x4XRjEkmwAVG7AZA
iQmwKiIDqZ5SgapG2SI/BUkeoo6RQp2uO/AcfKwtdxa0El5lSlubznKglXGQ5nGTRDHdxKYq/il2
bGNe4mtVN7uOPPBYwk1Nej09XnP1pooVJhH1sbHH6grCePpJ75yBi95Fk3tpBSOcB2O6n1lW6Pz1
qJ1yiin9FGbAdOIkc4pDnGspvd6qL6GljX66ZQedT0hxouHC9sSONWxiTmW1GI6GVjIFFeruHUDX
RUKIndznSKm6D9f8Ws8f1sxd5F0LzJJSMAGZMBeYsAIUawNGY2j4edrzpTnVDhl0sXxvq8W5b2bp
zSCHzu75TpOE1dE+phAU/QiubZWtKBH3U2Ivr2oLtV0QplJ+tGVlP2pwFjfxxjdwBbVimzFpaIHx
Xs6uRHaTIC152JYt7wDoULLygf25b/Ongcn9mg24IIC8pWpA+KXf3nnyqDCRUVrm9JKz2wdWkE8/
ku8RMcReU56WHaEaSm7ZBbZKRaPIwEOaXT3Ib345pF3Mhs/QymaPWviglW7S/61OIr65XkAUfBKU
4OdHY5dK1aJgGMnFVma3UW3L1dmyAzB1ezlnXMjophDI+Lp9U1MflE7EHZH+Kd93HDiBdRqQPo3i
mzr/hY2Z9KNT93v7VrR3lSqW3vieem3ohPGCEhYNjYzQvOqgeSqhg1fe6AeKT0FMRExRX2ZS4NS2
msX5I2vN5cnCtyKoAgsbNrftA4tbVGEj5DQhW+YStbwCUdnPHgjCfSlro0MUUcx7tQOoYGkDV+La
TPu95LAhJsdGmkVFYW9i7xrKcNdmmt8jLXTnfHZjhuZy0mdHfhpQlt0ryH5eb0zGiLK6jC+5Vo0T
saz00Gk7CEpC7c83Pknj3nag/iTKCUOz5/jC4BgekJMt6W4MoHcM3mTu69NsQ1yzfANvVFB7eB/8
AvadJBwQc4JwDN91pkHrr58KGl2sWDXmZ9q0cNADzBQw8v1Zfe0hs/M+IcCotQ4574ZfB+CARnr4
8sIFCt5wU1PIvpeDxevwVD/wVq0RcKqiG0dUI3qXsKeD7m1BwMbkTUoEueY7BOkANjTNHKFRluGz
D0ALjWTYrEGM5gaue5nC3wDka1FNGT8yhSxhGORdpd8UljKzL6wyvexd5MaL0V/RMYMA96EfgctF
urTtGTQR0vCXWMrWB1bsQdT0/do4KzY4cu2Zpwa6CjtiP0vGKyCVJ3YV5JRoEG5ERJln1NoQpEwi
wei2SeXJ1LLgdYI52sDFzywGWTkjOS3toYsDJGEzD+SDQ+sUGZGHDD1R1HNrJ97SleAG1NFeGwd3
vrcQnJXarBjzeycrAO/Zl8dknq5o0CmeWNRBtfMTFhcQklsg5XdbNFXJRKS1BO5y8ZcEPbX5qkNK
cwqmvF84g8oCgtvD46PCrXONSYfRWdnuVc34MECa5d+q99+yDqSxe9B58PIuAPP4dx6i/E2Etl8r
u8xi/DDHUiQ1aWSL+3JHxQmp82HosmwmSGTz81+IMKMyuSyrjRcnjxEVJpiyeEIcM1I/wmo7ondi
EdotEB5IapOEgNJbLPE5WjK+i8A5712XR8YMSfr3WyhVS3q/Q/K0usJ+ptRCf1X50U8VQ9MS+lra
mjlY+M8GP9BksZnLQMwtvOYt9ncdwLgRKqhoZbY3YMS+ujs60DtyLwMuWFQW985Jf6l8k1nvqzXx
3H2dBwAngpBz+QEkkVDHB1MXqJfDk5UK0r8JfW9JvmNKsFUtEgZkMurpmMC6cvuuvyvRXTM0yEjD
CuvP8sTwJKesBkPfD/SReBUgWSNzbsk95PFD2M5a7lg67nH1paFMXJ15FjxlytNDWpZBDPYcFu+r
VgcNIY2ZwmgxuFnyeliAEungzrs8MbYCnEQLhULA4FhAjtr+oVVbTuL3XdwbawpcBJFZpn1PtldZ
qHOZYjnZeGVO8jswFLIRePCtwox9KSleAflSO4Nus+Z0Gl027gx0CV2bvX6RTIuIL7YLMcSeuJbF
2k+qTNDB/Hiv+Z/FoylDMC70vjHgJf3NXgNLRe67/QRXmB2cw+QtnlHLhb7tLsEugXWg605VbHgU
voH69UT/oBHrzsX1wSCZr5zPqKTXkqYngtCoE3f6QQBew2jtJSb9VPkruVRUw7Qk7By646CHV90c
s6Kpf3EWShbhkAJX3m9p4knuS0LvfUggBClcHF/SgU/7gGamGXOedcSXAp8FnDT2UpJZ4I8VAjF4
KhRKj3VLgG06nDp8c1Lp875wKA7riQcHC7MutEOdSae6Uwc6V4VW8BO6AhRyJHhlbK5FjoWBO272
FHJBmn4x3s43Tidm3osIo0ZSoW+Kyyg48y+7VPQUmhTPfZ00E7idosNd7FgwI7bh0ebxfK98tQYa
XUQDLy1dZsGEIrFmR1K38kfCXmLkX0rGcdgrP/jwqQ2e9hpKr7GW6wQU8c7bOpjSXUCrLwldfDLx
zyfzswpivb3Sl+93JI2hp3f0rxIs+OFAK4r89m3zsz025YYPDizA9pwonyCuxZqyik8aXEww1GQK
p/0cmQQIhTZt/GHv7qjaTbMEDzDrQGhaVynuoF85gLlEXTnjstAbBIXOkln6oKYy1mWmNRLAn+m3
wPU3uUq0AliB1k5RP2LndZNCoAS1XB6A7j3dJBtCh9hXlA8OzmuK3GB9VwrN0DqlZS7PDni8Alxz
D/wk4+T6LKG4tI0RfkBOc3/aGm0wv/9H6BbXt3HWLBp2eXdECRy4CDBL8vD3ShkcU4BMblaoX07T
eh6ZfO2vsmpIfK+TCvS0dadi/btExvHmKw99cDysw1szrvZVgE7upYeR8iEXQE1PTrIs14Wtb/kn
Voe66desTG/SHR/k+hQm9B9Uav/KLYFRu9iLN2UrC8X/w/ngm+B344gDQgqUd0sG+AQhSI4oUxQX
GzjuY3jxvI63HiUgXRiebVIOo3piqjGwNXXjXSQxc5Nz4vjG+uC9a5WQJpLgXCv33u6biOjdYe+g
0Cr2vFLqQUikH2QQ105sDwIaY+kfxuckKUFegFzFOP4U1fiNBGvC4/+tbA8lrFFFN+jNM6Q7AQoZ
t6fr/CbO6+/nAFnVbPBsGxhbY9Gr1eJU2zR1kbQndB392b/ixzZ2WJWurxdF7Aj+jJg1FSz/WpAo
bY/zim6pmg74tkjKosXAvC3q5k9dJxDGG8OAkPAhBD+aIXbXCQrLKGyqI+76IW4AnQKhRXYSVUjX
2ewa8tUbCrW3ll8JdOAYDa2e1mC31OUDB+qtXEFAuBDCarhZe3Ki0ZZGG5XoXl31X+BqzfFjuVA9
mE7Cbm1XufbuVKQfpSeMgO7MqAYNZmFJzM22Ztm0Xf0MCsYCUCfFyTK7Nh+luxu5OEeUrsWx3vrE
zwCZDqvUQyXoWq8WrNWVErgOODWip55gf9jJp6hh47B/pPskwwBNKOCFr2GPvYTinatqwg2Uz4n+
Ohm3GSEmQovq2KQGKFaiMvJHlOoon+OafF3kCpyMkLRKbS1JYWGmWp2fvv/wLkej8qjODSwbcEeG
nODOFfp9gYvgBK2BSilpH4WS5NmmITGPIexWWnV8P+2h2vIyZWOgA8ooyy+MW6AHls97Hp7q6dJS
5BrJvBMZ9cPqQHvQ8H72GJ8gEFNrWp0oIJRkvmt9PDSY0MffJ9MWu2veCzt/ieeFo0uFFOX9QgCN
Kx/Xc7SySWLUIyIBLQs7mHFn/BEuMw6VqsbBlvAqSwVlSTGXypJ7CbQEtCE2cW7GgIvrFQ9qoLhX
KWlWD0K7GvSRZ/zzYahGKzXkwNVLlQgqJ+FgYngD2UHHptbVAQd6+xvDRx1mecvxWVdNhUdjDpfe
hP59GfV9TK9CG6ogQOjk5yqqSqJ/8q7mtuX4v2kx8heET8pUtVhoHs6WK3wDVgZVHAnBbvAFHNhX
jDylABndbm3bXlxZ4+xkmo/2tE1R0rAhmF3aiit3sK9YS8JQJGGyqbY+qDpquDUPecG2gqTB3kvc
hXTJ7zTuRK9oTr2h3ijLyLh7PkbzAxCYei3acztu0m81m7L4VUbdRHvrLZePmF3VNhSAhrH2ZjFi
xKsTmhw1/+4L2NuJMdiHA8LbDbGMOLqyVJ+n+wfTaOpB1C8+FSm2kTcVtRq/fUrprkl/lXdgzro8
jOnWTe1yKXfSFIX3RxcjIUszV+ECB8dKfcsaBJffcczB4AFLWt9NOzpmZklH386mcX6QlYiV6Hsj
oJSVFbSelNw49f5D6Rs8c9KqV6DV5T0x2c40M9CDGvXB/m98b+b/vdjqe/BaUG9M9TRK5+oiaTr+
FJAIBJYd1xCyNj/O6giMXZgZ+xSomK4yx5VCHojCg9A/ErteHP1v4ls8lMXTupQS3c8IhdPS8rj0
LJQrW4Zu/NHxX0uUBzb2ipU0gDznR2EN/TtZ4p6CVkJ8i6zVdj7udSXKy9mjyZ6/i7CzbSDMekiV
ot5+GkGQBoOMaB+kJ9rPKDOx7hLSWU2M+VGxZQGoSD2TH4y+A1bPjKym9eiDVUP5cARqeXS5AQYA
7eUAG2SJBsR2L4qbYX4NCaF1gY3EU9nB1TMOwH0AvK2RipryRpqwjQGvW+p9lyuotpqPAvvgf9cN
UsbZFNYBowHfaOJM1i2d9ApKTZlgUm05sh839bri17ADsAw0ljeTCIjX8cbBklky4okgrWLD9mYA
BOcMIOBG7AyT+YSFJa+Q5Wmby/M2MN7cnBdTlRbf7L8gK62+0e/mO1c550tFgmfkEq1xWE0kKRIP
ZShWiSff6E75ewbLVvmlr8pzijycrNsz/5kwtiEXfPYRgmzGVm76FpyfEx7zSW9n7FN7ML4Lk0hh
e9JyMIxOyD/UL0i/NM/+HVJYdgyw4tMjvDoLemhEgVWLjSzhmR2xRgnn5IMCm1chLwOd5KXZrhR5
9cBvc6IvUOJECFwhyCr6l62VZm1FaIdr5rokhR1L9FvRONA4qCH0AUW/HZP1jbbvs3oDTkIPyqee
kI47SpsCM9po9zsCi7120BxPGiAmh1VOBRAA80U/D/MKkt2biY077i0IuW+6mq5V85vK5zuT5wYd
HG2YjD7MimC8Wx/j7lFf8Eoy70m79VtUG+sqg9uR8w43KLmTlVpLsFL6b2Tf4YOKoNNl8r7RgyOS
7wkgwAP4iaLlj8WC17CZcoMbkp4Vm/x7IgK0HBgJnTqNZeaLREbQP3pMzRd8Qs8HWWspL/7hbZhd
Sp8guGjxjcPmE8FTsWsz/6WkfiYvZOeWDS/O7uX6diJSPn4te5K5SWG+SFido/NwdsFj10lXhaDO
/gmPMyHKE1i/NHSJR3sqLTUZ49iVydsxgJrwYUeUiKDsJSQbxI3v/D1IryoI7tDyfiUOMAzao4wm
ZxOb0ns4DPG7dk/rtFUmex2BTv4ebky5LaSjcspYeCX7YUDhI8T3kggAYV0/v1+7YZz20zCakvuR
HuJcUKXjWx+Riafq8NOnY1Jjlw/iGb/SgHRjS31Mm+LZPzv43SUcRskC8awF8sZv33nP4tY0/Eci
vmamxOFFMPdDw9ue+mHWwHui5fi3aABK7z3bgjAFGQS7auvqZkSLGj6u62xhTymip3+9Kvr7jxXc
aqjfW7Q+f7e5qT2WQfc3VGjSXysCZ0/vCuji7U7YjT5JzlNMrXNHmPTsESnyKGWBqCnS35Wy0Qgr
9KcOG2/nemSvSWuWgUG2+NG8cMqm508ZZxnffXGplwIE2B8GbNvOHiwIC+EHo7RKcROjeE5D9Kya
5ihtFG4hUVDEWyYFEfz2PKAT9ELIDS+bxPAUQKeXzpldeygYx6HkevL0KLjCt5QVnjLcSFvgW1L4
TeGnFurCKovlyaqv9B1xrmQ5++lCWZfdIwNPdYn/ElP1f1f3pouEPPFOkB9s83BSsZ5TzsqYnWIo
dKt2bdvQ4CBdc1Z3KsuJDRYVUyBBGbfenPxTAyfIra1IMZ1FqSvAYp+pUsEFszFjWT7/sfLNuIXd
Gk35zWDSFYfyCBpx2tT3L4Cri1ypItqjC/FRxjIz0D1gy29dZrcCP71fj2oweUT3wCUV/ukFiHx7
XZRleofyBvPptj6XSdq8i7JlVkgbFDR9UeTVqziAiqNQxEHb2LsOUzBOTPZfjKSuatbSmSpd2akH
aRjY0Wqcjln6On6VpTtUmB2WnKU54rcPruNZF5Ui5/UylPIChmZWw4Jy/pWIs1KMQtkX1PKpk6Nc
+T9nJHDRiqhiUAOAMmA7A/vIEd2YiYfUBgPU37nyp/JWlazRqOgds6DjUSxNRRmCC+DkyacMiDHK
sTVB8DsUzMG5kAvHifCE/Q8GZEM/h5Nt+3Ce6mSkv3w5cPSy6OGmpjTZgbgToewxrFjWNApweRyC
N0LHjShA30vnznRHBVlu5MF+jgT3DbcJHUyK7cPT9jYc5g/CzIDYDCoN+MRD3jhuzx554A8l9W3Z
M72yvDD/0hL4suc37hybHe9hvXHrpuYtM0mKdUxJy6l7pYm5akZO9WUASHqo/HVkPsgP0NPSH1Vk
FvQ5uEnspxhuJ3wD70VIHMgtycnip6OuyufDDvRMoCyxG6Z7CjUFnkzKFZ5tuHhnlRJixm+P4ak8
6bFteGHUpUYD5zMlJr61L2Mogjn7NgTw836HBov4tMrikvmknM7us4l6+C5gyUR/LzI/P4zy8fBp
YAEWMxqn1MA8aXSme7yWsRLK8jgu58rfTgvckD2LDNMMaGDWbTA/5jmitA6IoYSf0a1PK06Ed1tO
whhIySkuitTTBf6ZT7Ncxe1N02TM2aA4OF85UseMQtA6Uy9GC8PSAi7fic3SfGXcDnPVvq/YIWY8
Pj3GvPx4azbV7wzKnATa+PILoj6PgflG9PwgKqFNCgf6IzV89+CsGUUJACIO1jsMWfLNQ7YzfQKh
35aKOIywlGYdZM3dXe2OXig862gbUl4mdouBynSkXrsMddDEiN52/xjzYfckTCM/hCIqCugQOytc
n5lnnCbnRg8WAfjE7jBVyJVmO8/4oqXnUVG+ncnRnn7t7zTeN1qYs3BuKxO0fJDWfVucPb44ylJX
qgvHDwkPIkyYiyw2Oi1Ir6+PZZH8nhMAr98C0XQs5TGGjdsCeTvUqSov7bhTmc48fTHfba3334zA
dt/JjTpJK2gnANz8ZTniCG/3YSHNFjwOONq5djVRmbEIiDVRA2VfbO19s7yP2KLJQc6fyPLjfVRj
RMcRu+oywYTOPEDr266abRlfhMXt/ue4OEgNBw4FCZhJ3b1IiW7D5fpi9FE9I7IDFKp2Hn9SKcwg
jThjUmujbR8Pi8oFsp/PEFlX1onrJStOiIg30wzdhI5AX2Qmr2OccRN8oFKbubIeDowSogE8zOXE
HdYThfZjAY6qt5UzVEJ1ipw1pOnVlfMAiJzVPpjuEuzbTYLugHc9Q4Jtgj2IQbi9zAZxI1ZVoigf
5gFojU4ucPS6ETQ2tnayQUgz5SI2fYHv9rJuPwhXHdgWpMpJo3cnjGHGeXy2Xq3bPHeJpQU/s4K+
3gXzLqvPFo0cYTwGuynwX4VWrceTJmasfkUr+jTwP2oM8FslLeaEY28GAQhiS2EGNb9tTS7DIExD
Mbv3UUUeThITTynDo1BeIS0Z9zgwD6l/DAnOdzfJsaU0z3LFquJnFb9CE1lcppe1qIBGn8OYMgbS
1ASqc/V4YFM0HMlEG3+mRXlw0LUC11VeHXetI9axcSjZD/MueyVjg6kWSFL8Ma9dQMdRzzymDS75
BPmxrFY59sxcfpcV6Zep/kz/EOpuYWOk4kduEExCHUAhAzQV5b8TaBI8CLDUfoQYgZlTxJJhN0gP
WNzmhkzMG+j+xLlRcTOwwb0rY8sHfMcIFZRW1itYx+lxCeYgPupGu9mpa1Q8xPNWFKM49GcQdZk+
9C6qR79M320EqPtw3dESjakRHL1+god5LU1e2NXCo7KyPI97sxbZdo0DwM+1fzwJaeQVOrVtXNB1
aGgsZfbJpQp9QHGm50gMU7ZjrkosF94Kj/BxUSXZHhdglynoYLCDNNOEEHIkSyDuDhl3Zq/ZFR2a
bTEuiXazrweIuhI9GhuYOkoEjzDKQMpwG0L2zF6ujvmi5u4dtsVE40G8BGrWwrDachw37q3yp7Pc
xjIAh9sv2UBKHg+olTs9XK7Mu81PAnhDvMCHcBlQTPYFlOlCWrWaWCM01CYLHOc3ng85MNp0nAyF
/d3ZUOYW52dof3WlXiioU3bQ6vdVk4GdJ8KndeogI6gPLIPBrARGgpDUhOrSYC7Y/ttiFgUd4x2Q
Nf6FH01uHLsIoAY4WImNmrPJ+RYxlHySpWttvfRtpkwJxM+qniEIabyrJQr3OdOQ3DwcW1MsNgC+
LaRhrbIvNLM6XMElbQUW7MCPWAm6HSyeoGTqH6Q6hbJ+qEwFJ4m5byipCU/WKX9nMLDJXJ+mGC/1
yYDE5CYqKjUUJ1zA8dEZH4aBAzDERzL2+NZey2lqPX1GWESLGFjwpQP+Mb3kFWHojnba2+WGxEai
UdypPh8wwuTSkIW87IlzeVIQm2hr2JVY1gSPkQL/S38GFiQrNUM2WXPUZJXLntQETToEbqZW0vpx
QWCYvgoRdP1txHoyLsi5ZLCLCaiICMUbZGlOdTVI0DyZGE9Y6nXrKDal1ukOL7ViU+M3BSpT7S3s
308MVjz9pAviS3LU3x52OTbprqsCGWbIKD29P6PFj9O1JdX/556GhlSjUJLD++zGUUzDIkqxEnSm
dCtmbie+seidgCIo8vtYJCDJ9SRzhSoJQiHurEUR0pbh/RKdFFxgnj+UquY6zhfh88gr2E8HvOgc
Dooz6JJpTtAaqrnUYhtHQjuXiVVwENjm2cG34zrL22WXGbNbkQXOXGD96n7O3CWSV2T4HnqG1N+t
7Z9x0V8t4UU4WFSWzQwDrlt20Z6P8NN9QzyBdBsrSM/PVAHa3q0RArZxa7ays8wOkWE7irpmNY04
aBCuxVKIS9IVn5Hx8J7jzzOQSkVnIvY8i56GkGYyxiKiVC6Vq2hN1dMm9Ul+jcJrvVGMvmMEXrbY
Jrp1JSfpO5YCUtY2bzswSMApCh4NGTZeDU2CHSQFvGAGu61xigdCE9n5w6TnmelrNnS8TREs66de
5T1dRDcdycyLT+Uy0aWhNFGl8sKTAl3854vM7ZHSBXGg8i7rZ1HBnJIzjTX5IV6xBnoqJ8UHHZw1
YK06PmHlw0rIO9i10rpa2dukqqu2xR1gJlU5YuOOw6KLosI2ctpR3TjBJJ5Z5/nnTm1oRrzzjkIa
DI62w8+oU7BetYKkgi86eCW8xzAVLB34RcN1HjbAq+WA5jLFvGSjnopNwgFtLRjg9dFjYnvsqf3l
mXrCmVytweJkXKjpwa11sdvT1XAlbh/3gEi6LBPL1n6Ar1vbfu8yYXJVAUs59SS56tnU95D8+Qqa
rmOO8oyek/6wHc7DKlrYX5Ehx9zDlo5zTr+F3Wt45AD8mAfdwrbm/CBScFSmBcltvXEedI8IEGnE
joK6bPv28cnzAdTENbscVuDyleEHqcunLaN577s7KEmfW6pXfXOrYhzIHn1Lkc3YNTc8NgwbI07V
rdjmd5qj7rTiM3p5f8jXteoRUUuBzJSW2zB7u/xCVtOPd9RES+pDdae6Gcns0yf/tTqL7h7meDEn
0eCgqwZzcb/RwYIQNFJm7qlexMXUoEzFJTLmRD7Bur+GoCw9Wt3+B8f4VKFulC51zcZVOu2PXnL8
j5dANdzrWQqKLeOHRyFnBKknFYa2gQ2ez5xy4sE5Mrn72yM4keYBoxMqJ+APjjqiwYV3vVx7Gq6R
9gsL2tcRMF9SID/nU9vsKmJEJiIaeFFNikVnao+jdjIFpjSLGqVjljD0TWU1rT9Ge4ur1kLdjyWt
hP7rIIHeZwQjO3IZcvgc1IExfzjbwd3YEKGsBsqYEI9LuscfwnR4XD5S0HoAmeU7vEwpIZ6v6B0W
MeOB0d+AL6gE8Hx+fnN8OmFU9SgVv2jusLJ6D2h5N8bqg24g90CkN1W3UawIwplgZY4M8VOUQ3nH
Zy3dI5jCiNeZ6SK7C/5OPVRPsGJhdhvk1PLWUFR0KzP1Y93PQZTYwDizFzNHWoYE7cn/dBl1jYBa
lok3NJIdQt5nVOFcLeLE+IIjbUuaOzmh6ipX4kl4r2f9m4/FOhjzm11/HYZO+GtvzljACoyGAVFZ
jWMfD1MTAedTnHEZ0SQoX0f+mWgLI+B2G0IeaTLTQCV4zX6VG+hqUSHMVbsfPuxpj3ViY/5zDpED
t5gqYsBJPq0JPLfpFqKBZVRYFSjwi9yLJpVqUx8GsduppJSxJp4i7C4dfht4tJNmnvwhPsUadsuh
h28wX/phF/bo89d4JVqbMkr2LH03Qq1+8Ue+Qoklwq1P9ySpMIBCoiqIcPCnXaYkhU2YMAzOPTDb
+P4Tfpx4yjjdhX4anYYCXQ7HHNQfMbqN99dhErVrb7mlyKu7qhrFUvwfMkP3bhLG4vrHm85hBjjA
EcS7hbg5rtGcoIxBnPulJfw9XLqDRvp+rcar+LIjHwaFlr6qLlhDYllsAwXn3yvcVtYR3mN3vXJ1
g+HDYMSJpUWkLUTLB3x7OK/Bxr8zlu62+zmWehuIL/8VphO0yWKC4I2FV2Oklg14zO7AaaTlT+op
vbXWSs6RGXtgvn/nCKoxTuEYus8QdCTB04cAppZDFw1CwVAe7E/xGCYk4CTn8s/EFhmDBG6fDLFe
q92hGjphq8MUamFzPxCoa11jtjjjeT/UrfbWfXbKrp3QhSh7v+JqmyKjWtG62dGZUD9Y6rzJwi4/
fuj039v+QQBuU7YY6QX1j3faGofhAu89bvQyENHG37J2shuHz4WKTsU46x3Jr4Gfm7KhPDO51id5
INafj8GpWL8lNx18mICgtE3/5O/L75wRZQn/ehKhfyF750zmnSP474nbtPmR2NpLKZz/McnmP9t8
ZE4nvZFAFkoo3CBqllHZqi8P02YM4UW+1DKe3dbiF6/N8rS2BsOXEb/BdzUECL38WkNzPaRh+Exk
Ui/ytgsErTOqTSuz/8WEC+dW9V63e5MAbKCBNVhXqySdvVyYP9LyAe8hYDRwL/kWw7gYn+uYIIsq
HyhGR4USbVTvjkqv5bonu6Wk5zs4uObAHztn56/hJ0pPktjNJX3dkTUKIKtIQCEaJbo/E7cjWa6x
dEGd887U9aiWZuY1JNDlH5BF2GvaTebCmBwfA5zPggtGwcRjyEMtAAOszE7HqY2SS+I2xHwX4NN8
u/yzxBN9CNUn3ldd3VFdJCxaSsrmHczr8LsQo32cN7VPLT3zDNnautUzD4NJu517SB4F5AGmT4oE
YPfJS5VX1akLAzxOY1e4ROVnsk5tL/xHIHxSHlxypxUl6l13d+L2nut+iOkLeb0cPk0SqPksmxIj
En/IkYySS9+S+bfba65zOmCuYRVaUcRS6Y8o5HlNF8mFDIqlJmc3qwbziAabf46syvVkQT8XSRwj
8SKKAlhZ9ADTSCDiM8y9Jy7sVaXJM3stSTPPuJiTtM2ATHJ2eL41TpVwgnQv5leznMUKloQdiKSu
xOQUdTP5ljIMBTTCroP8hlZ3LwVLYcfFVmzMSby3qQXf3tNKX5iMk1PmzzqvIwgL1g+DHzFaaW/y
bC0IwUE63CGv4PBcMzNfUWziGe2hSSp3CPoLIyXWk4NUrYRFUo1cY6rI8gjB8ALARnyrksXLvOr/
+84CM2clQ2FM2iVfXufouSEl5VTmxKR05678ryb7Q2oHaFWKvWKPL7207MpxSXOGkbN3PbPbQDkK
K3yJpR6olOkvGlPdj39vMczdq5w8z4r1zVM8dXUGKiogiEJOF34ThBQN4drdh3ORVceatSGQtL1G
uZZGBar/ky2elTxR9KbmQ4z3YeW5aFl+/vARQnprPfG7Ct0R+FnZhvS7yEII1/JX+2nbMETlG4Sz
aqVXimoJ/R/m+rz5F9SfDzkcy2S6w1msUEwwYzsdTSVFLYKpGCCLApOGw2lmsIuLpHNU1BBJ6B2Y
TudXYy/6wfCvZwKML5IHs4D2duW9isCV5flM+i+bf6bIqGJ8X9NFSmu71MVyDUrhHoiplKaGBLMB
bFURD2qQozwmBuwl3QiMjoJrgGmdR2rosP5bTEBu856a4KslSIxYzKMDeItlYsz1yFemXqnwTC7I
zYs8cdboriYV4ecu28yqdtOiBVhpdqoWTqslWVZVIUq7D6INbWQkLuE9sXsShn9UK/6jN66ziXhG
7qojqYghYVYNgKZ3bgz79yytOoBtpFcE430CV8k0F+EUj02425WMFkSKmvvEu/0DCRGucRwvmT+X
71jC24eLsAyxg/jqTzrMYNuR/7wTWyZI6J0vmHXvrOuISfUmALWc3HgFRlSrrxryYS8StoGw2V8O
xgD2/ogD2Yhw8t7gx2alStWGLvXsjf6bYHucuy7S5rkWMuiDchABYfzyQCh5Rh9qgnvydfxHY4vS
4xGrZbuOcBloV7PhjHVm8lBda0bU6yl6yUuPgq1mZZpSLI4Z8n/7lpO7YqaBmiHQjfnn8cryy+jC
ea3cd1P4xSpWjLp+dXuAo2nKscdWDFt1OKQd6Mo/GBUATwL2of5KGXgLb83mIuauqsjAfmyfTh96
EQLGGcTFzZxAbmN9RXTRsxSF5cCVi+uytN/D9f+vsxGzGvnP9TgGSLI2Bt7TwBwU/nX3jp3/TsbH
S6D0Gw5wtgCBEnwKMAZCAns2bqxq1JIIs6Z9Ht27/JV0Uu+wCIiKoWz+U+NmjrZwbHOTiNwBc6Qz
Uk2nC3OWfi4n1bkpSaeXvE2hM2YS1AVfCddSpi7KL1hxGp/3qTBNnhWx0RITukmeNbTUPwBPGtzd
RQfoHw8evNGV1pNl71dQXojbMZCrjFroWUWWHlM9H4XrPTifyTsyTBekrxBHiIl5hgGDNhzOTu/K
iKHo27P8uNNx1HenoqLr2rifdjWiHIOWHX8ohxPgBgQcrR3yt817Wzp6hesJ084q01+EjylNdybI
bazAE3nLQz95KQahodnW498i6XHRTAOZuiFyzulHuxAFXVOH9KdtsjSYYB5RqrH1MCLgsi7HWoK1
RryskEzZyfcfxEIlXBLzQOVhpwczo//8mnWC85F788Dg4fXA5cPOCd0sgysPsaYmM5G2q2X1qIQd
dLXc4h5yIVpoDxcY7xwO6ioyFhUMhBM3Uoc95Ev2LSzLLnVGTk2zv3V+Hh6sLbLtMc+vT5pN0w4n
XLy+U2uE1rYbfkiqs/pjSw1ekPzPLRoUVV2Rw+eRzBC1PIKbD7sRMzP6BQr/ajtmh4BT2TwogRuH
gkpxliPR0I2nwxVmrTWpZWp/wt5hqadSgYdF2xRXj67SurobvFLmj3GzsdcaNZFMpNQYlyMnRadN
yq5hHMbW9ub9GE8d8g5pxceNYa1WJtrJrY5tyuulXEn60Nyk6WTRmtQz5E+stoJFjzrttKwswFo1
Dh6Iac6dWvbdjblO4OklmbxG0md8zPGNMEYlyT5EhmBgG8HNBwAuRGqMJ5/6p4ufAtHBns42spH5
ZgaMV2GBs6Tn/uijwqW93U3vTd+kErnmFw9OdubpI/oKcGuMBo2QAZhVch51WYvpAvi4qhHrnLoh
dRPMYztpzM8+vDSmF39ujNAIOTYj4psIr9s2wxC6iGdC8kXA8k1mTcKfYrR+7iqM4h7rzct8KsKq
i9S/sRF8KASa85u/nzopLKxH6l7FsFRLrRtyyJ/+ZdNvo+j9Pqk2nJWxZ9CYMgApeqWkf3OK2Enk
bYsZfaF8LvyEHmMKrMUkHaVhIpXumdQhS4lacSjO4lMwBg9xDjAddpbKBK+0aHyN0uDrFvSidO2/
grzVjmbvKCVkuAekTKmsGvL43JEjFOnJ/jOui9bX+uuDTW6X9DHqTLGzVSAHrZqKw7MYilGnbMV3
EOujwU72KUPep/C8htgHIEqBFugIuXdSnpbKfd+3CKYy/m2IdxWQavOxwpjKwoF/ea0xaIvqSBB0
ZfyCv0jlqhKzH5ZjcpZw5kKYyx0S9goWIflFqa93dgYJijdtbaTeumiEysvDLd4+pJtkS4xHScMa
zLN9T326x5mO65+EO8F4bpp7ZhsF1UkkEJtokT/fwOrwQTynca92SbUq0yfZMjBkNgnswjKKHheL
2RHy6uj3C6ddPdAmJVrLLTe9dBRq+5d+Cua618FxwCjk4633f4sYcAeojLExUs3RO+JRoK5Cpj0M
dybo60sp/OrXkHLSivd5cz2GkNAZCmDY4q3fYZBzPb3QMeEfDL/3AxFcxQ/MqrcVfGFgFt7hY6qt
7ZQaj3LOAsXs8s22UMGUq3Y6FmfPq9ay2L79D1goa9pELODMpexFyeNP4l1kV8/tBr2APn119oJI
OyOtJeq73WWKoDN/wQa6eUAE6g76mZhnsVUHw+faZWPAcF/2NKSAr6f16ig7hZGV2zChS8s+uque
aRCmCaMQ1wyMJ+3gH3IgJkSuqqKBRwNJfnNnw7Vdf7QuIgWuEdocAMio+LrS+jwHi7FOWH82n8gt
wtInd51UdLvnnEkIu4cfCqZl74ITVgSl9WUsZjQYlQXUNCEdXMscWAQera2e9JEuJbzUqZI0l5NS
tb/hClXRqg9dH4sxG6Fkr7A32fDPeyvQL0FA8H8JRUAcAs8HpnLl31oyI1qUDk1mFW0wLui2UaY+
bZfjkeBKPc1lgzIpyd9lJjuwg0hKFGD9BL6Tlvy1rmlniUHiiTIUtttTBY0dXeL20hkiU5QyEj+o
tcULvMTAIJyG8hKKKScc0H7d66uVQB01RKRvzeWHnI+7QPcVSJJkOQ0GDu2vJ5aqE7Fv6J8+Rr2y
l9kcrB4H8Lbc+en8t/Zk2IWBhMNpUNLQyOICP1CgbtMnOpFpacHVZ39zJyzzQvP0l1ZFm4YmEg/n
NJKiZyTex1WlAX9h1HGk2q47sIENQSSigyi6p/nEQoP3cEQA3W7a/dJ907e1rhlt8x4V/pbyEn5e
obY50wCvyNgNlFKK3axCGndoOaGF380Cm4j7JEpGuwxn3kLwiL7aWNf3aXi2tiT5yQjHLdD/FHcj
fKQqYCD6b/lf067IPJQatynt/lmXpgtwtnm35KCjGdySdFrYlJfLk35dz4DehhUfLBXNyjSJHAKE
ScPfTJ78HHTncIfrpX7QtGy/5NayKQd19SkFI8PY8/QGsd/Az+joZhOYrPHXqKwpJVjioEz+YTTJ
5w/qJjDhsn42R99nwoAyEG4VRkj2NqIKCy7v5Ymk+D2JseuR9qBywXq9IrFN4jnuaya4Esu6XArT
lpTSAQZzm6sUDUnffRKDD7QMGjubz0bNpNwmCpSOkhc3RygagoWS1qi7xS4n79bNGAJWzsRfTtng
8ruAuNsKxyfKw+vQwQ1FgHgGa9Nvpc0t1cFyqkb72AvNaYKiOkh+kwU5vUcb8OUzSQMZtC6nzTfY
oF6+uZUlIXiw+Zg3fPQqzeppysdqGDDeVIMt3g7Blr6XWjLGb3sHhbzY/m2YPU8hW/L/aDRh+5qe
A1WA35E9DVEXs3RGQAcAbCkPZ91CdGmiz73LcCK0lbpiKlG2O7Zydv0eYvePyv62ituGFseCCuKF
oJpak68BUsRqR2YNhh16r0dC/xtDovxzomXWjJWSHhGss7j06RStty5WE8h5N/901LmPynrjiVcp
RWaoCeVr8c3NYjZAAZ7CIFJrsWMYa8pD7tBqvhl3wt2fq5CgfzjQZQ/2/31Yiepno0pcdPIr4lDV
vU+dtyAjFCG4AlaqyAD/KlOF7a1ypvDBAkNjsXWvj6H1zrZffEGYncJ/YdvhY+KXOHixAZPx4JQM
1Yuqj/BOhgQtigtH1cNL9xokDCDLqXahhvqGEAG6jbAV6Xv8cTCfvdQ4HbaDMJHi48/pZpt6S/vY
lpV8VG3j4/WazetYBv7a53uPaBe2I/vobrp6WDdpURc3euzo/8botBgD/rofYSYtZIBu+URk1WjF
dhtE06i63Rd0gy59QTAvoo+LnCI2qR6odR/c0Ehm7g9JRpg7spDfoxm2skvccmB+8Ac3shvr49vK
F0ZFXcuwp4oeJ3CIQixOeSCCMPy43PsglXhYkZdfVxI9cr8ERuJukWd1WwPUNNrEjLSiAV9D+YyU
bc6lkyStqSi+at+imLg4A9bTVvoaHV6jKl/XVro9AJG/CyahhZMJDsvTMS2T0KYWZY3oFnnt6JbK
uTCSw/pX3ABepo8O4DKmAoLp6b5CdqqE5UAW7SQy+Ht24E4h7vAbgfUpVKhOv63fsJD/CKmyF72j
VktobRdKpmeo5UASRajnk5QmqB+AGGO2s1/8lo35jcq7LUhtc3Or04M9y+nRaEAAeV82HImi8nZS
lrvKOspdkkDqNK75K1kpvqQdnYmZCXXz1kBVbSu3pNxs0pBWwtcXeVnFnhS4CIw5S+0vmkhBFoyV
CjXZT8VC36Iq51qU2j+SRa5v+qTQK0NJHgnCMLiNX2xV7KXYa6nvLjw7vwPPOq9ZHGu+rsrVN4S+
7mjtFFmhHuI55BhuEgq84CTxis3Lk2Gj+tY4nKDdnZcAUa0pu50rq/UgyrLDSTC+N4mdkaiI3fMU
/BaKVOYWsCcRklc2ZqnHjkMg3x+zc7l0SOfjRnfoW15cNmBGUclpVktcZHCOAWqmJg4AQrD3bXEH
bAmfuSIJ/hWBGyp3WGn3UhEjiUZUPJ6OXmdKWL4uxpZiROKbLhGslH+oEXG4nHvMjgFNYijwYZdD
v673pO1MoxPzJzdv4bME2zglqN25RTrztAkxLMP1MBH4k0MI/yPdLiJLokHjUIPdfBr++udNNJyt
WXghi1MWIBCKuta4qTpHI98Cm33akm+f/1q3KdnESIrFaX5Re9uRsoaNyWbkHhxj/05MD1lPWF6A
qpWRtRLEdSJkHhYidfpgQ1YKpmKUJrWx0EkCiQtgcdsflj53Y1AE7Wwk0G1uptk/CYaSx16x0UA4
3KRpJ9rXWscr/dVpRNLZda84c1fJSF8lPGQ2sBhU+EfsGxED2WQfdCZ4kQPR1wbXrCCT/M0Gs3AA
IayIybbmTel+eX25wjzXHKAuxJum9Xz1RxWPDcOWpFTBVeFOx2wunS/47DixXGA34V27MX3bzF5o
SX7W1N5n4yJogo9e7aAXXetIiZEImpXnk0c/wkK+XfiGJqYrko5tBQjFf77rFqlEWqqND0szOYMg
VtMy/SCd8wyrXJKetprqcZYOKQ7MTyjv4cltgRomQ0RZk9Trvb9Wbkd4SOSpOtUteQ5QEE/XoQd+
ObfVn49VOlJdrkSot8+YDJd4cKWGshipmxyZ5uz0a42+fDRixZQN/AGCWf3ZVWQhLPpB5kZs1mJ6
4v+WaJDqgcM+eKbs+sEqQM/hf5ACOoqKuxtRzq4V3bE62wZwNFK2nGbJpTnD1lat5a4Ss0W3j5Q8
n6tXmvJRKsC8a0M/kVFseC1r4yrX07zlSqNnJYQq+Izhd3QRrPgL7PZet6GGqKEPH+t1u8dqL3Dv
eAWoqkjjRt1/sI58PD89bBI25QRXjaUKPw3mUkdmGGgujYZyJ7bps3GDBPQzFmBzDs3R+sbfUoMS
bGwDSajU0crtJ9Mc/h5IbbthMAZ+L3w/+n/TN908/HrEjRpMbayBDg58gsuoGsY6JDUrwPMrgbyb
v0dhxOw8IxDBy8u3Td9zWiVOviFDUXSevdyrvqgs33JPueIQ4F4dftFNVCPhi5owR4hFGMVnICsX
pYWmKnm8gIxE0PBwvCV8RiI/waxhetKBtZ+Fb/iiqaDVSHGAiqFrWo9vC/NZI2WrLYXzIp6mp9eh
ilxaAfbhAqi3chD+QUxqY2avoHZU5WjEB4erRL4vcCVixV5QQ8BWzinO/FfT22/2r8iVDVCSeKPM
VnbtGuOV6NnbTSi1y0T3glo7Wvsp8M3lImg4v4id9jJNFxnO50Jqg2Xp4fHSYxbesTaDdSMx7yM+
Dda/0HdAs0NP735rpt4Dyf7ZOttZADGvpMi10FPPb69rNmgMyKtZCGOAlSQmmAhX3DugHw6eFbGc
6PXjtYy3oxWDi7DUOpoFuLa/wjzFHhITL4ASfO4ZaUJCfQ+cs6DS+RMFTwAyCzD5VVcHQR3ok4g4
kGt52aFoP9nAc3apIP3vHKw+aFE/XmkmJO3cAH7bLN/V9bKn/W+geQ1Sxm6CM0mio3Tfr+tp5UF5
GSe4b2/yRXa6S0rysJu+doIlWZYMbEqhuQAryDZs1ah/QDvTHoXHKk1WRWsxyM3jEIs9WC+A8Bfx
pyJNLYLtjJof9qqs9XeOdFpDPG0oOrI/w1TFFWQItgVr6xfYL570e//c9T1f5n5ImPSor8rSntOy
7R1YWvpfUqZvT0dK/TMwlDd1PnQAY1zQ6qg05uE/S6y6dR5+Ji5LnefplSsDZHyUBCBQb+2kyxMU
70rssG8jndmNGyNtoGPPZzyeG0uG990t7Pny8R6UiQoMRaepWQC2guaZEuANv+K2lwG3MBmdbpzR
35QS/+QMis/JKg166DkFNt+gRlA5yNzcLyBm+ORGw8deFIgwD/ejpK6dVOpL+6yzYBayrMCkbIi8
DBqrdjw4s/lp2HHvS4EpMw9G0GMd0rN4BLodvrrjGIalMCIILWp5WBDouLigLMvFVi1e9SUqV9ik
QkBKS7C3/3fv9KZDAROeIWj40QrFMeyMjrw1rOK505L/g3F52SO2BuNtz5Zcfmhm+KrzslMtvASh
psbKYLDgGGnoDeI8CnBLWzpyorVj1KOB8H8cAl3V7P34G/vQiNWp87V8I1kGqx5hZ3viICNEXQXC
hVTK6HUP22Od5/gey+QVrRDB/CGgsQt9H8QgKYuNcu1g1dit/dLs7BaWSbqnjP5EkxunzEQTF1R8
La74Wy3OJ35k1t/cFntaxZ7xnXtlhYFKnhQD8FCvIzdpVoNx8mxbFxuQqk7FdJlpnslbog2+cEmX
VuDyoD4jvhdzX2xaY6JpNxAfNtsFV6XUKcAvelqdjgXT8k6bOdytsGQ+mOLRFL2xA6TjL5WPP4pg
dsNTMVh+TI4pvGzAULGzEJ5TmEOf+Wn1JCLGcmHOFvv2pzH3+d8R5cNxRaxexrJKdYKY3dO1yoIe
r/dCC0jh5zjZtei1giji3VXZI7fVRK9t+0R9OEXpgrg4y1BZmv3Tj/x/lGhC3kCI4khXdvjNXHm9
law5uYRA4WochToPt0JgvUWHGkH31Iqg7EB+rqlpb+h0XInwhSYvyxHSRqK1q9sS1xauZPO7pZEW
VQC4j29V22gq/X67x4S++NOQDOTQDzmBqYDghoWeiPPAnZsh2dzBsGXFO27DcYrb4TO9YZpQxNL/
I6sssHiVEpnoOH5ki5/Dr9As5v0ZBzQNkrrXFSq7N8jjLmEpI7W7hqGxlIoi6a27qe9SogyCAzyT
faYhmZ9LJ0cAWJjlKTmu9aM2VOSZ3vx7F28AxWllvk5k5llupVyKQIQQ5IAeohK/4Mmjk94noeRY
HQ9WU+hcCaciHW8UXsZeRNYu4W+6yVeb1oQC2LSNZgZaE86Y/ndt4xoX5SOjHVO8+97HEEOL1wNb
/ai+t/q+TE2/qKyoab489J4wgy2+RIm8IXJ3yZlqSmko6AV3BrvR5FZ5aZs2tVblgqfbIUKb/Ajd
WodDnUA4P9E0OLzL0f6y+xebvqJtdAwm4GTtCiAuGDX4dyte7oJMU6WAKyHQLVgyLN3WvG1D52vI
C0Mbbfk55quU16sCMuLTSLFuOzrNtLjPgROxD/zZyIgH6o1cbqrxajZdvpfPdKl+D4ede+gC/3kX
BesdOR+0pJ/IZ91kpeLj5I1vOq0HnlX9fKD/07zJX7FdoLlhARMarx/mw9IjbIF8Bpnq0IZrNEAb
rN6ceEgtGF5eUSLr7/bXOqX+IuH4Uw9E8BhkHrWu88BvvYxlbtyvTqcz/19mFPmDHscbJ40OzWDK
a4b2dtIsLqALJQ3iDGHzcwQ2TOOc0PMmLwj+jvHNl3FFmhDr1HGfHKAyxCtTv1dTzBytth4HmIsL
zBpv36XpSxEFg1RBkGRwj5ZWCPBJa/aCxLStrCEzE3mI0p2IibF5JCHmgwkJswBKUnW+NHioX6rr
NkkXeO07gw+BJz9Ji+iD/j2MR1exzecRHE8mxcPyRV9b7auHcuq8cj2nzAJllR1VH44vzbzWaI/M
w/b+cc6S9JzM5dGzbt8DLXKX+XT1C8ncf3bmEgtSjsO8RugR12DwsxF9k/Ku2hblBi/pXRPBMkLN
QCf6RZQa/Ez6lsrZTGy6w7o2SlbnxOlCFRroxhPpHJ92iLXNbXT/GSoFAtrGuyDhQy714GopDjaT
T23yLDZ6qaU+vrWggCu5irb48Qw6/VLc1NkSpGhOtMaxG8gbgNjFhHtidFdGJVDrkeG5hL0h54fm
O5HqxxGVzQ5dGBRiSasKyYb8sBqz0w4BpUIl/z1CmcM3Lu724K/btOSGIfsoL+6kIhLpG+hHzylL
scxu+JYBmHfetIfaBzvt1xTpY9w7JHQdT6+2nMQu1/lkEd82S6dyTZfPulJzU7yxJgcYLXximNzQ
dx/9OsyOMeTDAXxg+YUE8bTCn/kyyRc2WKFlQD720F2JOBspeN1mths1TpowAHU4stI0n6ibCc+Z
nJyBWhkSeTIqkbeMhCzwhfRXRgCJR8a+SQMg2XRwqkHUPrLiPscJ0p2Ssxf2vGkpTRGf64ZZozT0
iKAdWvUuFgW4SUFZOHCdKvG/df2mQP1CwiLkXNcZipN95Ig979sH6j3tBdFl+yK6yGu2/rA+S27I
57Ttfv8SjECsyxzI8SkTrbB4bkvXfOCewAQ7nWMgXELSP4E7104MZsQ2fLJbHxiiBpEVrOijkXWZ
pZ10MD7NbFMfg+lwtwE1NpxwwR742fgwEYbQjDMxEqdU8HeGOapdx3RlNcJbwfUvEIyyRHk/hT6h
3/qcw9vozfZ0LKdHNelhfA6rupgr7pr0mogzuZdXGUIUtP/u87AFw6X9gZrKFAuRKVt2snRNIJwB
vru4KBNaeRDmLu2brckjYCxADIEkPkEFKLJMAS5JlYwOssgv4PZagsZ4X8JoOL+LblNJgxzfVNMn
3kb/+xYFglYRpq0pFVY2slKcKP/NwI1L6BTpVYGCA/pyqJUbakY0ljDfInCDsHkw27jNtjRJ+D81
cWwCIdAUGnOhQF9kj4GElA8dtN+MSW9uu2NF5hZTB94ostCXHJUKJ/eZP6yVHvimEHpM0wOtUE71
hqGO7RmpDOMDAmPvzONnmk6wSi6BIIcTZYSnSpsnrIF3SoJen6DnZzGkZRLsRX17Q0QSoN1wA8t1
goSYnGUXpF6OCzyWiVJsSqQQ6FNVhcJ2l1G6Z495jiD61XzVA56B/EINZhUWEH/nhuF6y6Ao19G7
z/DVMjxi+PV16atU3b2RKcSwOOSYVfb+KZz9xgQfqBDqw2SPcJxuBsWq7QWM8rpuWa9Ps71irs6/
J6Bh3fXs99yRQ2Q3UwKxU6SZHb9wE2kFAYEm/WflXU0HQ0vu1EXbVrC/Y5kmko7hPuVDxDSM4qS2
ZdAzD9i7Tj5d/rajTlEe5aEHi1Djq+DdEEWnQJUALNtdJkkmRozKBvRUePXds1FhIp00CBwLyNnR
PzAbgsKyVKiARNKiy7ehlZC2YPEYHwnj78Xv0VtDIvhXDhHSicvEvrkdlnwovhK4eiBIyG1BYTAc
KpNPzbhlHXe70az2F07G6icDQk1fF4z9lsIQEKFZf4i8Qys5SxPpoouliGEEbvoGK8faKcTmwOg7
eUTA1fogyokDi72aDGkul9g91kzi1204MYJxpnnwn0tPmWhi6vvznKnrxp8e7bgkvzLJY/2JdaS8
NnWhdrLyaNypvbqKezKJHsu5+ShVFA9W3BJxNzUFXKPgOKI1n1GxkMthTu0E026pESPvBSIWmAag
NfGh63eUussNymEQ48h7NBs7c9WgA57A75Ca072RQz4j5ELG5uEDdNgNxyZNkjbF0Hux9gCDdUV+
QQT1p4oCQTGw25y1q7iosG0uSDzyyDeVFeS+MOQJoD0P9Huc7UKDr5xrRwx1mSztkZHVzYbizkSR
Mkc8V4E4d0a06VDWypVLhBzlrik2z0sD+PVikNb9Th7FaSAs4lnWwtS7xrAldwgh/TcqQ8JiaxTq
ADGcLdpHZYr38p8axeAnyWcQuvDjdA8Hlxv+4re/zbYBiztfNpoVTnZJRSGJW2u1lACAr/StfF04
9vbRSD8wWlq0Idx8gKNrD7O5Q7zZWzeFJg8rSIchrFN4MCmp+bDnidpH7theIUwAilDpkHRdORll
4GNZ3nngbsjKd9fj1+/7zsKqxX+HqPatOkAoBMRESjRG85s7de4XqXlxt8m6vLmEPnYhzz1PiFzu
433p5t0SfROQa4kQjLGovk2VelMfyz1t4OgoGbgEU+Aarv74dEbEUEDEfwDCUSDMx9MiI2+v/WEl
lPpAZBxjJ2G4uYOdjs/l6e/gEeyQaqkROr3yyux1CkVmANEHaPc/NKJ3SLUenmsvzBsWCD/KPW9b
2rUkr039VrRjsN7pKMYXEqDwqiS2rbBi7MxR8kcTdcUKlbYhyDQTemOA8dU1aDMnnLEBhIF+5FZo
64MJfxzHYhUMMmReCGFcdWeXr5o9OqOCHuM4SHC0P3wlLc5v6MvWyqZKbKiBEQ23Q5NXVjtIDIFI
OKgt5WKY40Oyt/Dkz4sPth4iFWs/0Xf5mo+EIN4A9Rbj/D4l5SBpIhjoAT3JEOr1txu17KDkVFkr
3RtDS4HOKwDoWPDHW4APb6F5bm/ir7lucNnXxtbaDfupIIKflmwVKmM2qGbVZEDUuA8YQz45pxtW
KFapqA/Q9R23kGL3xt24tFzsvquklCqOhHasjmyztYPQAfzpvx+2HnLCvQxQ23oGPACtqAgTcMAe
g0A8U5zE6Ep1573apHRdcgOCKpmAspC/AJf8gPK12PlcLu7A0Or7z84Iq5PtMDz4BKzQG23vEw1Y
jB/dMTVbE00YG326czURvn+4IdOkxFnCAGc92hL8oelS1F2JkZPx7xmK+xTqQvjL2GAvPRaeEZXc
X0Gk3d1cATlCj+HsEUJY7RZL2yE/5nwTp98A385cdHQwKY8WMrEi5stW0cgaoI5gmqHvapa0FDXV
N8erZhWuBj+qnQg5sostpGQBOn78S8Mo1EDUcW179xWDhnIUR4+XA1DxY925kDXQmCgwOtw/OzGW
VajOnhn5rjDS1WPZTi9HSPqDBlefb/7Ue51tylZpR8q8xptOiN76MInwkFMdksTCiMsxzzrqcYm3
C8nn0Vyq/jyJTLyCrHCR6IR5SG7G/EfvP62r6G7YKb3EKGO9uPnJWhRapF5SVvmLUzMbYTpMURul
kpqp2+2aPRCifLhM9vdMF+clQ4OXdc+4EgVl1o+80FYS9V4f8wioBV/MKdGePgNTbKAXpAqHwtUD
AKns6xU5seNPus8EnK1v+vQBJ+t8qJtjL3nDlpcfHIT9c+BvTRVBq+HwG7h5Z/2ilzpOTQFWLwbQ
zuHl2FQ8D9w70dCSQHHj6Do37sTnGIuYZfccvpsIeOZifw5Dv5IBvq3BrKJZqj1QBOUnLhO0bowE
BuiDDFWdCiWhq0RX1ATHiVKPKLrS6o3FoNlCMAkSdHQBP5x5FhoTKz/unOM9ZvvCcCOWewMdz2gV
9QgLn7UjG206WvBc3jxU75srN1wXGvfq/1l1jGh3czA1xjgKt8FCxA/3u1Seza7iCggyQ84MMvcX
IIN0cT3DFRKbIdZBclNp4c5Fl3Xumc/ZR2TFDM+7wh5gqyR40Zg9kXLH+SO27mHzkE/QsFr25WuS
w5gnt+06uAgb88wAtxmvtwBkKpMS0vJG4a8iqGoZsS2TtxzephmQIRXJ78igEVMPeZCcp5ySPwRS
f6DmQfU23SYLxB+u4RuZ50kShQIMD9vtnKlXfdIlJd71qtjjdPtPGZch58NM+V0iNDu61v1/sop5
scHS1vdHu5j/RT8rzrHzF3NPU9+PzPtPQIyUnjKznQoJeuAO7lvRKyC7Uv+7lwBjpNE5bkXuEQ2N
hy1C3ZRIa3J9xliF/QfUIpRGjbMTst3Zwi61NtVbLwjt4i3R1DCs6ELmPFnkCTTO92LT1vJLH1aS
gBoA0jEZU1o3CtTr3vDkq+HUelCAnYcsy+zg/vHOw+DU76+REUQtOidgxQXudhvI011DuW3miwZ9
I8NycIPyrkagwjdt8lAxis7hDVGkzp0Y1xsepk7pFRtMzppy+pn77tm0f75iNhUDztVZ0XI6+Px8
ejMMQpDSupijHWNj4MQlcYv2AFlYYPs1akD5cE1RWJbD/iUcIyG5JtfhDI8oxZOUlweWq3j9iptU
lXUo7tqpvaevKPRUHFAlOj8xFyvWjJhKM93QBqfS3dpoqUFuFZAGV4bc9VpOAjWZUusn7/xxP4o/
/YlkZIan1Grnxf86uEVpl8EtxR43jgmm2Al7b6UMD4kD78ko0AXJ3ppJIiayiktu1izbdfmtXoyH
Tgcf5L3V1yoV2SLVvWUvgeRWkhGDv8klN0V7TNBCQJij54lrUzCpFGiHMOghKsnOYnpbI60DlYkH
FSMQ0zK4PrAoRd0nAEgUrEHaXAyhuY9BjTPKeb8fRVxxnrpYwJ7Y7AUR25Gzrqd9JgV/fqwHLbnu
4flPfAbT8VeCvDPDMwY8KhXc5FiNM68aIEB1j2YZykCzbfWmJpSdOPAMHwHCdi0XEdX83D9QF/40
nXtxYo9S9HEIODhEkAl4BWt9U5jRrtMtChnlsONohlKvGdZRRpAFjnAy3eRNlTeJlVJlqwlAzFcV
ZoX1ysb/EKVvGjeNWvKk+Yf1fg3yeKRgxej+9Dp3UlwGivgicc/EfrVY9tdB0X6Hj2DhOob2VsyC
rjqZa+3isyKF1cLSPCFC6eZYcvtdp62VUMQka/WO4K08d+Nyl3QucQqUIeJPWW/O4hU9xmCAT30k
t9BPKqeowBvDBmmBwA6Msm1NzB+p7T/EaKcFI8iJ6n5Oxn20/2G5WvhG8Utgdk3vt3DMiwRTO4ag
c7PU1yXMBEti9+A0UPM3drp6Fchgzs8A13CtEvJd9c1ix/bgx9k7jrph133/x2jQLdaFgUqgNu6R
Gs2WWx+EWom5haoeAh63dx01QcRkTm4znK0BZvghzZzMqdzBhv4e2gxiRC9kGcP1fKDdXHSSPfw2
JkyF1O7ZNy9EHaoXHh5cCGbg/C+LSB7JVSoNoH+TyNUQ0XusKWlU1nVEMuwio6fdI2VUfl7mbYcx
z0+WHIUK+qO08dA5zFtcswk7O6ANoS6R+qJW6TNN1euDMleq2Wx/a1teAwRl1VJ5OM0W4te7hXET
swf1aKJxHeh0piZ9j1e1iZXLkiNgbdLN7w0trWUswuX8TPhyaOv97ZYBy4jZpFmI2WVxUC5aTbew
79kvHZRpkFyU58YJ6fFhzQYke4TYql1nDcoSzcIfBjfepby4pqgcNi5u6n9rv64UZUACJWWWg7qB
A8S4slIEf9bvm1NP4ZeO+x08S4nBls35oV/hCvfJUfhUexJzUQu26Eh0Cdm6l+4uP3pY8VnPiUnq
tJcjVLTJ3FGs7u3ywvVX2m1EhYU5VO9eK1Enva69MLbsv3GVx+Z95TWE2pJcPZsS0DcHpCl3Ps1M
NRp4LJEG6Qd3xG1YST9JK2kYz4CTcD8gi0TpoBDQXsnt6hDlxmnvGqLyuDVnwi3DAQLi5YBxL1aD
eaqDpD4aA/lNWZEnBvnbEX5a1iUvBokFXCf0pySGxvzdSRbQBgiPRXDI/wc8LwGdAqaEV/ixxnIp
Oew9kNDOS9TNY5k7wQ/9jbSFddb/ewaLws0gaLbupGbejhKUqA82N90nl8Mnf6nyc3+mZFpwpM2w
ETvrHbMIJgIjKg0xcnbxb0DROBVKHlE1VstSpN4RDvklKJMsZqy5x08ywOl+HzJ4g9XGyC/8bP3E
mL77WvWomFv6ByWygBDHsptrn02q792+ZO4rtEnp+g+KhGXiGYujMNtAYxN8YzyJ8uDEqGBZ8CJi
aVef7u+tI8cmDBFFQeIPp2Or9r6SeuPIzsDrHklxR3MfHaalLqyFI5T68MubFbWIRxqmmBlIgGGs
/lef2STd+mKjOseviKdHBbm0ypZZoSXBitjOYay4l2k3LaLsEK29gIF7ys+qsdTZh3Hlsf3B0eC8
ZoKcf/NIncDQDBT48PpFJbbh5aHBnTbkUO1l3p5YHcUkjd48+4dckFW4fleX5pkbXg1pR8UZ69fz
kxTIDYuTnnYKsOubqdeT6/RSVWiwm5SCfHjj3Kf68L9/cp7IT0dRYqE+BZWMxtheh/dpyYVIPADf
NPNXyrDe8iuCD4CbJkK6zL4tXqqTBsCij4wwOFQ47Vm6qnGBAKsQj7d7yXTbwXcnGQkFef5kKlil
4iwWz1Bss7zJa9xmANZ7HXeU5iyh3+Q9mEhQWf/bMHzR0NTNvniCBlygsLE8tT4XK4iQpK3t5Jb6
9HYYDzvt0NcUw4rPPUb7IDYH+9Dfz3sJmXkQp5ZMn2mLMC8dqfmFdxHGvpYYcwG/OOnynHRvGlhg
rbIc10eshyfwpAlJnBls8ck9NQpr5A9fNz3dtHuibt35ze5TkrGIafkRAR3f+HkOvS4xgRC8qC3E
s0z879sxmgoZJ58WgmL1cE47EsllCP7s9DadOc/pgwOtiMdP+2XVTrNslAKdSqTsdSE9S8ygzxH2
Cln2MbAemdttqsQ5ilmInM7ehcdghP6bZ9Whyc3rk8OVT1HtuqOMXzGBQUif1ExwvcbNLR1vsPxZ
CQsyC4rwDC8ih9n8VsFq0Q/C53PONKUsmIRQNhLGTjnUApGFeCfON/Y7NMmiWRyWZReMN5VeOyB7
rUmHS5ajALuU+DOSBhTL348w5nrwTGf+KQgbwg6K82KLFUM/UCTMwbw6i9bo3QbDB6P8t6OFGt6k
h8BlXpKiEGlPCGfXxq6k/FZ9jLiWbG4DKNp70WXZaq4G83Muai6wZGTgD+UJd1U9xCG0gOZ8xJkG
ORFjknBGHv5qPWu0tDvi7Onp/q8D10wsSo+LtYKepkbLgWvUdSzYhXE+xkb+GyIVtK+EkVbt/tiL
0jn8WQAKZKnOjgxl55vsklAoAhOmrN1K4Hdj8zRXzBLQeM4sZFgFcZoL+Q+XV2yJRAveSgeGzmnr
6laCSgLxyZdWNtwd41UAmLI68rAsL2M8r7NRumNcKd3TWULM4RD5pU1nhawpmPfzNRofVXY0qsXj
dObPVLlfihpIdIsnKjYm4STIZPHx0Zlz4KTmBJQA9JIHBJyhYi7gTcUZKHVZqrs9+EI/p+0Q+WA3
Nlm5erfEKKrCFyrd+UsshstiaM6mmpT6kXCrRBpItyP5iVZ+f9Rv4oBq8dKXSKsz+/ynU5QiVTD+
eQ/4xU+bBBkD3Os+vFf7C4EaRY4hNgnSKD5yGjgaF1gkU/ZXxA0g/vyv3asthSJVfjQ14ZintRye
dMt7r9g6IGYBGHMOxJTTprBLZzX6aXJFdxyy2l3B8VYTpKoQOfC6CmNLX1QDJ5ihSQeQ4BEFOuTC
/LNC+t3eCAEoRAmABRiPjNya7hFeWxx3K/4eQrOHYD5OMUh2Ss34xXeY8POXWgkwJgo8Q/OL84X4
WXP9ysw1VlNMvObbPFf8Jz8HV873LbO8ru31b9v2FYHSQGPD+Wq9C9YHzV4Vb+tQd+mqcnw+7s6P
62htTG6MDfJJ+JE9OPOCUHcxBPI+Aq/aq75ROVMio1vFG6wz9kdwZnsuaJB+kdhNR6yS8jz48fDM
ZwXwD/HWDLFWONbtcXrYDWHCgGn/teL0Hsv6arx/HPwjNsqEdl82fHRBrE4xOV8jE/M83Cp5iZRy
I3CvY/YnyWTdyzor3IWqG1rA9BSJWFNiKHo5Tdlp+GKdUgMbncAY+x8JeCEGnBX1lcZZYZ1aTP/L
j+qUzR+VpVjaXAZ/z8LPRT0tlo20qfUxCawVOccOYvk5MJjh+QUyUw/h/19nPvyyMp8S7ojoApWh
MkyLpgJ+JUHcp0jJvQzPSPDYNJCrkt180VKxESGwjyjKyGj64ptcJuR7CtZ32Lrj4bde4nBaMMBM
4LhSCEFoKr1s3ZpWp6kE0MK9tjatDDFUhiVyhUQOAe6sL/2ZOF9TzQJCOoXSorEn8kTXfCTk+yk6
QEySaYl+QjupJzJuXEHRk1/QvrNCiwnjGmixlu2KbGIDRmFHA5oZDM9ROByeELNIaJMVGG4uw62R
1guTzAPSpzKUpqFOZEvEAJtVKV+XKV/KsXNhwrLWv5h7BSKdMHKUSxsdTr4wJNssLGz+5Yv8qZ3S
LSOo6bfgu7eOt1MMGL74mNYOxgb2YFamgQKu2ev864YWGoKTyFjslK/SYN4S2U7/nnp5CNfO3GZS
L+YyPwhVHs7Oe6ulj7Xajxy/1GKmWIP1FDvAU0dS2W8uWIXfq3vJy343f+Y3cM2Ha1sVo7w2TzI8
nIJQrYs1l0n0xj+hWJr+D/u0RCJbJTFc//4NECHCye/amT9RcQpKJlYS4+iaYBUwzvszjsNXwt7d
t+5z2kecAUH8bWfp2eW7+gs5W82dODIEO+jP4etMaVXGjBob8dAjaONL1IJ98d+tm3/MllvyrFdH
kWYpRPO15AQYh6+iuMZlzQpRZeBNdjO9UCLyQSESiuif+g13Hdvynl6ofSvz3O11wuF9KDxBVVui
p6ownOCIRh3E/1W3PfFP6BnFUyXgWCIXF1F49Erdsb0TQLcDt1CsRsoaqxF89iBJpMMsSIwh/EwB
f1pLip51gSlEah0tmy4TrIHc9gJDNR6Kc1iOmWpUtRv621DmApQBE8WePVYOgaY2n+WQVoh8tsoa
aHpn6ATPwejMIlaS4IvgHIyCDf1OOCQ4rJxFsX1ZFypIaKawQqS87mwZrvWHD+JeDMS4Acq/PDFz
PDk0/l/0NDs3w1jDEUekqODQYjdh4N5BJCAId4DLQpgmPbdd0vtlI1CehGWuMckZBeJmrHFuBHib
+4ZwWwZN9ltJxw5+2wyOMbXGdnaHCvuwmDnnB92L2i/IgMaC0lzgDL2tKbUH8x1xGM3/leK04Lti
iSbqH0F5VwYYkriq9xk6D7XBNs6y9S9PRWWR6ZuqiNnP4G3yndbMIXl8611wXARmPNvDSs68vHqU
nY4+PM+1z9EVhu5LGcyj3nQgG2of0P13T22pgDDbFBjeXrRZJaU16rSritJIm6ddXH9lQc5rZqhu
NdW/CcGgs3LCrVD2DgyQpaq6MsOK+0cLvuIgNEkSRYJv/gbQ1BTYZ0YbHYMzxC0xrYl7uHWSpFys
4ucBfehLIiptN0Npd7YbGHxj+SRsPmwNZ0zJV7+s9bHVMns2wOeiYeRoodYJ6iGieauYGidPZJOu
nC1at3Ov61zg9nASSl7RGLxxgxFSG4sPaMf+ksMI5qOsCkEl+v73srqVVqFCTc1QOhbeQog4gjIa
ra9Wy7scvaQyUIBV144Yb9EanAoK7XmmQEyBlZx8K31JNxutR8sJNqKKvXsyt3i+bRB9u0OW02Xq
Ji9kw7d1l1t/9EJb78Nf2PKwW20iDaJ1QP72yBoFr2QMn4HPl0rvSWROCj9pdbJI69Cx5NUbwDa3
tJnAG2cM//6wybtqT4fdt2mbwG+scZgKNj8Z8949HtgRlUnRHmHtLSO0zDjkBTHbsVbcjxj1HqmW
/wWKebd24/scEtVpAaMH4eeGycH7OYpYg3Sa+sFVlMvpzS+jNJhcwYthprBqSsEadb69fZsCoyUe
zVFbN6yDEcxn576mXZaVo4e7UYlhmoNEulFubsojZpHxu98CJ9zE7hnOxwv1WuWbaTPr438dC6Wg
5Br9MnO7dzCZTNlz1pkc5n2OSyCIFXiiBtSBuxZZHRAxydOHX1Z3o5HpT20c/9GGb8kEekwGciTY
doaQ+xQHYwujrJ1udyDbuEZ6QaGL8b8quGYmCSirVPbapGDqJ3dm8zXaT3uaH6OgDhDTZUIXRjbe
9C82KIGSqCGuoNi7aLQyvWh/82pCS+sCXmwA2AWyZmw8EU/Kfm0fGPvqFpGIQDTRNcQacOUJF/8D
pz1t4N7lVfEHMtdO3aLN+WVf8RToRvryHw2GmXRODjQNsye5aCXCQf9AQNJmh51RV/Ity0W76NjU
Q4dkomn5l7mPeNpRswm6ozhQj2IL+6AfOAvCAm0oHK0NdLxIPENAqidlJ11UGTTBZAplxelhhsuR
GYGqRAJQn9izvrkoDM4q5RHzKdTJx5xzXdF2NiSAPjH5GEwmC4GZZk4/tl7LLjnLKB1JrhS1hkcy
+4ntlgU4apXuM/6wIUmyL29h1+fTf2ugJiev8W0jRmNIbw0xfFRoZHPAjsv7zbru95woyzvd/W6T
OPHasd5SHLK6mQtxFxKmuaWgd7OUEt4J9RUAhz62sAhc4BKb7SXQACw0vfULS9slhWYWBTAgdpM2
CFs0AQumlQAiZkT+FuFICbY2MJDunEQXHQ6bSYzdxHVKAbv6PaHyNWgL62puZVx6Zz7OgnFJ7cpH
W35lrh1d7CRUy0ZYkhmmr1a8oTR4htRUJlhX0JGPikuFxS8hubjnoVVYI5IhozBx+ZR4fwDWIZJy
cj2Po57EtrhKE78x44MBkvycNE/kcqOs6EmQEzwMugsWGKaN0oWzKQsu063OaqJmTorZcWImqFq7
diOIDcXjzKYYoGziGEyQnqMvF1p2pk2HkUw+Q4HHV7bT0YmiC9wb8WZu8Y9AdMfEYJvFAz3MkHi6
NCL/SuzbcSmseBg3mVHrvs/ovz0Vmsze38IpkR5uKd+HO3RLNI31hS1RBUe++NwytMvkZVhv30ox
b9Tx7M0HhwZMBuq6Y5/aycaNvfvJq5JoDEMzU2eNDuQyj4s09Zf+0/MJ43KofHwFeEeeL8BmOexg
aHxcGOiB1YMgBa5nJbuCAXKLgK19vBLk0IffIY21eZvkYUvJ/JNuCCQW35wJM8QshKx2WsiuG5Fh
rX5VZcVgT8W1MmoqRy5mfMweeq30/hIwmbu58OxrJjDxUpbgkll7dkSixpUCT8hvWg4bQUQC/X53
067VxUZ2E8U1lV0aPG1+U39x4byluoyhyQY8C/zHb1tgYcQieW/KT2zmQilGTy7HY+8iLqN/LINc
mwMKJE3z0TDvO2MdUSDU+fV5BDbbmWBocjU8attqjjIItrNDSEhLy1pc9NYiWYwcmvgR1SImFGBE
41iIgHb0u5seAFh5IZmFR3kNFbxpHJi1en2+hRmOWAqUQHTcvz8c3FTY7RT36JvqUUb6+OERyKqh
ynVuMlRHpBLezZ0sxvY8x0P8udItC5voc6paAICMJpIbiUhmoomZNw/OU1PlBGpYK+VO0rDteoxB
A1z9GIevL6zViK7YE53F323ZJ1LIcdlkl8AzXdEL5R0psGKQA6dWdXFImJc2tuy9RJSIdT3bbKsx
gyqfzljPiMnvF7o8J/+59+oLWeKKPt7R+HWbDSX7lCxqXAl8BljKUXBlGiDXKOe0JwchOEI4mzgU
FNvkpZ/FUcJBqk+BN9xGPVeHTjCwh2AlaS/sNER/ZhfvWpW2sV1J5NflTyOCD90ZVDPcCxQydrtP
YNsJcN4TnvilgNNDXKaW1BuwlUffR4NhqXPdxdi3oF/VwNiv8Y0X4p/F78CJEKfXKIrAZCGnWjuJ
F55r6PZhGxl27CLPhaxJqdFbgItDAJ9EQ8mzs2s1D90hKyQLewoQ1e/TTQ3Xa/5pRAWpDjruM/rV
or09W/lEkcXVT/+E5K1lPu6HTEu89HMNDoPgfW3GweFTVHpgzxV61mB/CNiYqfPaB2vU1Az6c6yd
P2ID1PFeDONy4HJc++OxYDGUu7NjTkOwBXD79B/nO7MNhooUx9n5UfO8gucXKBo+roTjas2XjM4t
HNgqCqgu99OX//0LlD6N2L+7sYfJQEQ6X/Dxvg3WsdwPYKoC+JTKEZz1fAe2Ff/QuSZsqnwP0ylT
8h9SVd+eITqhQp7RicsIJt/gY2Pmt1GdkGwWnhm9uLok1vK0qmAFBB5uNU8Gs7ljm6OIAVA0G7wR
x5khqrWx1cZAg1uvUr435J8uf0+W84iN+1XDTDou99XdDEQ7bV20m9t3p/CWzjGo4M08Qk9TxZ/2
dQJdA33FTqpY9TKjspl+E1GBFuT3vZCEXvm+O8QkqvjdegTll0d6q/paUa/707uRptrKmcQQbl1H
Ijk+UH7NpAJdqZmUpsTNbMiwRvv2urHrZieUYxK9S+sjahFk8MFbcVHlxsRiEqE38Cw3ADVk9gu4
lq3EwIkPnoeIvyy5/lCHIhpSmsVjAC+AaZs+aWkWPTAumaE0ME+rImGzhUATnRypdUaL+XC2Id0r
IttWG4iYgi+nQfJbC5rKBrKR+yLokkoKF1b8meVVzMnVB2xkgCiYgwtd1XOisluXaiJGOEiRT9ib
89YIL7gmTjDa7th0R1btxJCfaUOA4NeNIC5x0ATarHCipXxsvCKrIxpE/h1Wm7kWXcr1MJ0VmXFR
vQ7qFIb7f0f1sahcdW1ZM2AJOCUIpDUyf5GsN85lYVf0fPDaJCtwaRlGUd9D7aHK14G+IyuI/Ai9
0rbUTUnNst3vjhkaVWmn9zkf6O4/ZvserXMJz7mGfgaZEa7Ru7+vV22tQTTCw9ZpDF8DQBUCqHQS
7Vr+b08uxkminI7TIfFDai0Y+S7uSLymX0zVTilhcGj3Sz30I1Vt3ZyzW11g9CmQkhG6wwRUzT/g
eD2fTBtLYaBRWoBQhCqFbFeccXSK2nhpt+RTBSR1U1w9roHmm6WVY9klLEt7+4q/ZbIJI9CgyoT5
7rS0oJcWfvMRMdgdy+Xnp10VYoWmploWkTPMP56mkB3Q893YW18kwv49rQUebh80Haztch+AWKaP
XPLn3hgX5b9i6Z5va0C91ax1QGiTKX/M4ixzXZIEBThr8oIk5WMlRDRlPKTb0u6B5UH4gMwKIGNo
6wuyPH4X+evaVhw9ymAspqacf/gbVKh7+xyHKWGaY7VF6JX9YDAFxRm95T/b+hpRDlGK+8CKtHh8
e8RBEeJi3QmghBliMjW7gxNh+RePU+KCQYVqRi4vgJwqEUd9Wp8I1kvL9ZyyGDK/G+T5qP6v3YA7
Uqgrs5O8uGqC4hioGCXRkOpN6cnvoJsXyL14OLONv4H2dPWzvmzAsQiAiBBGKcuN3AhLr6y795VS
t/5iW+RiJqBIJbgpbwK3WB8PeCD/Htwasx3omaxVQfwD81djxukDbRB/UvhJklYnaQvnO7oKOUot
iUZcN/T70ouv2TYUILjfXQS6EgXNyzO6m/Cqe6aOikaT1jGfXWGCrUotUPhRmYsc2MTzab/oH2P5
KpkP1Stsgo4rxGHYuRuC9vNCMckuPHJGD1EOkAhgwhlBWEwGSNtkLHtcfh8brgK3U5Kjh5rJ4sgB
Qpa392lVv+O3p2xwORsRu+9uxEkufLj6+j5+C3Hh9abViExCtjm3PL+htkEIYQsTDsLCIWSTbXX/
OkR6rlra432C9/p/wqv3A5w4OQHAZcV8xNOP1KyRznalkw8r5pf3Iyae0GSSldPRCt7G4UC/2zv0
bEuryG1wLXOie2YyHTzEPt9PzsU0Hk9bFNy2W8xhS8UIWWDyxJv9OBI+IkqBffSyXWfdb/Qs7/Vt
GZBsvVcflvsHKXKz6TDPpyDPpJQSZTmqRovXuITx4c/RNhR4DdunG89XtYbTBNpHtxo9rXUOs10S
eddiRuY6BeBjQBMTY8Fm5CFl+TA9oFaYmE5mMdeeoa2ZoVPKssHilMibqKDvUBRkwH+c45U4anan
brKWaa+oG5ELkUER7ygopPjveuEE6/pkeluUb+EMOCsriCjSlZ+6+uH6JhKYsCF0xGdVuUFhapOa
cwSOidToXIsbHFP+WkbN3yen7++nQYL5ssm+jXnrwJJZlaAyqWRtT5EXIylcA6l4njG+td7KK3bi
89Cdb5Pmv+FJmVSB8SR7uyM9fYAYEbTcAS5RHsLMI0FQdYEeyuDDxNrE7ohjPKI4NVfV0txlfgbR
KYRZB10QxNTWASJhXaZ5yTj9QjG8z0x8AMmVYUKwaev47lJ+ywMjP1MjoG4F+y9rQ4F8jz5RkTpD
KRVkNRPPPAyiA9Ge/4tVPljLobanx18xTNwZtzrc26IftC070OcqWdTX9zLqREiP4pvt45Drp1T+
XCyuVP971eGeizwjmr7ZOgkcy8tz5QhQYuQtqkuOVjQl5DPXgj50J59jBk3vM6GwDFCoQ0vVUQxV
U+0Q0GbxGe3niVz93A401VTNPUgadFDdiceBVJLYjry+9avT+zwagSzG4ZbO6kfFttAEPoLFcxJq
3i1ngCPvW1cioj/gS/e3r7iiIw526XnftdeCqhgHzoIOwqG7iOkWYLGUR56Fb/o2YsQNGpLCuZHW
fe9slI+tuWzPytg9woqKnYmWBDdReLG09vmLsW2bT3Hk2aHq2m19WqstY6jnE4omA99Xvg9MOg2C
AnwGBoRyT4vLyv8l9nU4RRLYGqTDHR025d0/7WK3UAF6pEAj4PcIfLii79pqXsjxDkTHf0uSr8Lq
mO46pYcHHfnMCfdtgyUIOW/BlibIm1DpKaRftV+jVJW1Oe6aa4uy52uAdEGv1ghf0ZRCgmwmTBj7
Jo2iqRRBj5DvtyD0g5d+oaJ9oRPoelKaqgA6GzmRJE2wOcvYr8+J3qI7yr9uBtlLFZUiKsoWpYiF
RMmblKq9o79PvBy6um34mh1+htRkcugRjZsMsgesqTDoYIJF5Qm1xC7I+c0nKxiqwMec2LeGY8hR
gSn3omgUksWBdnXcI4gCE/ZY5ot4j/QA/lP+Z710RXuvmsCBvRmHn5AjZqfRc4bsG5Xy6JThE5zr
dIF6hsPjeS6ZGxK0L57ywnevmaiK/0B5mwEPeHSyG7sZ014KPgLoteYRHMf3rhAUQIsCgck5TgyU
ywqybqVFHB5/auJqyQEeBCPWPcBq6D5moaK5zk0p49vo/83R6Xnvt9V0IaLDSAN3eyqPw/QPT/X9
UyoLfoyeztR2EdghTGywVGniGopNtzfBYxQ71DagXh6j+l6nn8Hr746b242dVpOlTWalXsCyD550
9o3/RCXukT4IFsPLUMcR79WvoCipADx3dYhQ5/Ou2+hHwsnrAB+6ic28I8o1GXi8VvbvrQ6nkLP6
W2/+yBUj/rGVnZU3uO7cFYdnVCpEPnIp8X32a76UZMcUhi6xPWRNp6TqSlZBiWUqXtly656gdm3+
dafoGLF1OvoqUEpMaqKXIrJDtlE03V8YV5lxlHCEEcQej5XRtJrL9DTA1yb3bQxIcyOj9l9gZLT3
nYGNf9erV3khJIJnneBMDf+sKj6P7J1z4egWb6g3jlS5/KEYqeezed8dXL+znwXOn2irQZKpPmNr
aBx6PpnxR0cbV2lj+pTsIUxYvYLFoxsCMfzItDT62NGDptXE6jfZ5/k7E73j5vE+idmY4kP9SIMx
KIE4SVniy8LaE+SemmJ45ObSUOHhiAjBzwugGe/fz6vMNEE0mm8oJpqaLUYEQDXvGmogdAw2vjYX
TB6U3MCcrVcGKvZZI06U/5cq9FcKUoiaH6zObRQsLO3hku8iCZtr1aMIccH/jnzkR/4LKlktURiL
16i5dCki7rqivpUt6+Ohk91mLFyg9xXnXMpauIr4wvA9Kq06HM++T118oxHog1Tz8gClGkzemv3+
2cosb+s8Q9fpbSBG4pWxAaPyIK1fSPVrwxV4OmpfG0dhIlI1azYJCU7EE+OTio3xTsM/NxRywh+j
yTts1s5/6sTPR4UYil4y4oQSO4FG/jaPd9VUbBQc/flYK4Ymon9DE7zYKtwCbJqhYSW08yyRbgQj
iAvniLqpCiBi10kh846caTrbedxQjGs3IF1sZg0xyI1D/83alugg19dv4ON8rb564ZVvgXzcz6xc
XvZHH/Z+eDQzP/kud9qifuCaX9mVHJ8KIunZF0TODnc0/djNghsMLeLTl1dBXKZYaK3ZU+mYzhry
9QEcz+ZRB9/bJwjob5h3TXJ5Jhtqyh6bBC55ey3jjdaO6M5DXzRiUgE3tBff6a9iGyQsr6AKyAeu
Wd2yZQDV5fI73x8QYFCHxgoYReq+cJCm1gHweXKeekrjmLDMnLXDVyHxxLcHwHfZNxdFs7AXY3/4
GZFzglGD1cKHXKKfmnerl54NqESVqWdzsiYLL9Hu8bu4Y84IFuOlWr3jnCKQ0/JJX/DBfMhcwwRv
q/YaeMQMA9wek2C88eGcoDi3E1xDHCKzUBHxWWmryybflvK2rGwDbUJl8nFHFu0WzthDakLTxq3z
dKPMT2SSMHub5fDRuSiPbwJLEuWgGIKwfwFg4tabECQyGUYWTiuNmDdCsjKAAEOE7+kiD3T9O3Hj
3lFGuyMZ3TA2iGcUhzBkAiviagiIuyPsdua/se2wFeR7CMSCM6GpCNXRyj7CYtRouwJrf0kcUDFC
i1koWTbe+MFkOXAqid5uGOf5wLxVuygY+0nSzZQ8RlY9FKH1VpWkVt7YqjtiZGezV+iE6y7+T2GK
8FVh+dxIlhkfD7Xwt8KcVlZhTqo6CfeXTlIWr67E++kPy4to8uhL9O4WjJs/5vaHAzFpf+agtZ3r
ibu0dzzSA7huQsuOMIK/uHSvpu47nzI1ffEOqeLH9hR1x9a3Oqelra0uuOXE5JooJTA52P8RNF8S
8h4i9Gg8EOZMuJIpEpLwCAwuxWMexfGlKY+fN+ckpqpin3yGT5fCxrYKBt3z5SANSx51cZTIR3nH
abHzoaqsrNBvEYsThLvF65rc3Fre1sd8U/4KZ0xS2y8O3aUmyYBac9mx9p0dzKdKHcAamtgxj3s5
Goo2HVOUWCI+WklTPYmbMN0H8AK0V7k7HtfTDN5yrH3LyUs05F2VG2O09deTsXlEBAxOysqSgv8y
G47QIu+RqFcnXu3MPmleCLJ4wp1544zM7mmFoMuwrM6XqQ0QT58mAKduVLAJC5mXEoy8oNPstQi9
8BvvnsOyjwhNodkA4+4nLudWbWHZHSP+jP4NearfmOImY2t6C0a3VTA9NpCETIdTrhdEjnLQgunP
RBgPjOuX0JSDg2d/uiEWf7Gaphd3hKv8dxnbeto3Lear/G2tPUbodsX7g81owWaeE2dcAQyx5g0w
YWER0xbykPA/7VZ+ZSowcfKEY8IlFFAsF5l1wD590bsC1crHO4R9sfS1kBmny8pcsIaPxabGtONK
G8EI5mkkJdK1fsaaNiR4biBS0wSy5ZIjsaCziAIRjihQhMXFyVNB607FEMPI61S1GcLosNw3W3Xl
An2nXu5FBPRtp141flTL5Ik9BYEYnl9mjtqEa1xKInSlrRFZ8BLGS8jOl7nGqHmBJRpAksWaV8cj
0mj7g1ZDJOU+9eURyBb20pZJdkZIlFsuNwJqMgfcmjsW3cH88msjCRYyI4vkxo68f/GZjCotl4rm
+FsJYj4zCL9+Nky+3DJF6L1nP/HtoXtHYuMgr3q/IB56jvSUzLP0jSyThG96mTItlAQ9ljW8WJ05
L0HkrDlMS3Q+VNvVv8WIOpe9f11IwVKvhRvXys421cwwZyG2ke5iWluN9itGYx60PK3SQzfZ8HCt
LrFcNtWmSd599QTXHPV3MoyAR3L64GW5+ANH98DFzc3WvQOYCAjFcVHbQeNqLIL5makdrlEqnmpC
oIonPguEiZBiWeSgHM4KMguKSvSU8mtQg4rfXdNw0m7U4BovRFo7n4M8MYf4dPu/rGvgWk0DqL6q
UkA2h429zLrSh95Kr1kyD/zwyYnNNflnaMCu5fABsOump8jO+MP9NmdHvEtStMMNeYWFx9Hc4RsY
IQpFvULGTEed0abnRScIuCZS1iyVk239FM22NDLclejvbZ2xX9KnjIMxZFRSjiba4sC85ZGIjV44
2fIpnt5yyHOne4F/OLyVbe0WWNLWTKn5kg2jgXEe1Ftby1cHtOmtcNc9HX1s/LEk9X0UgbTYIPch
pY5BrC8hQL9+qp89RZAnZM/OABtm4aY54ieH5YQkSWeJSWsbaUufWa8mF/bbgv6Kh7AhEt+nkur6
kK7d0YRLx8tpXC0aw3V9j8Ce0lp5bdOJLIr9NW65sDd61NNLoRv5XZOwVBbfqbBRVp8ftTe2HA/L
lENZcDJbP2bSpe+ow3FauZ/kJB0ssWJhiNtWpH/s83q+EHgmDCc4r6M4x4ebTHDI6m/WQlCLsSnQ
eRLuob2UzxM8j+k+c1CZ3qKw7EQZAXOWwF/Gdn2Y0BINaR/kkBBhhO5eG7ANoZQx33H+r+raNKSY
cqBysBl692BG1FfdQ7nXd1nJHQC1vxWuVwgKfrwYmxxnVyuAdHWMpJj94udfdPOFB21gCJiGg7wt
vtnTt5+9Z0fuwJobkyJKai6siqqwIYanRZUlJSm+LPtUD1Hebtnc7hB0xaOEi0UmoqmxaN8NnVyF
Xv73XTyWtCn485EaOcc8Sy2X3xVSueLLLiHkkErt6QCLbVCigs1IJxQ3qoyGXxJuXOXAXli4zzl6
zJqfGSASSf/Z7GDIrjVcruxzoiM5Q7CE82wpSa1Ay2Zkga/CYGiU0iMWvKocALgnTmqWRW4j+HRy
BX0/c4UGhzQApwINowVUUr31Ka1EEWcZUyDWy8WjXn+A89St0+ueb6LY6snvQc/fdNLWArjPkliw
UBDG0UefsMXFoXKbt8Y+qUtpQ6fnVuicm+PcQzOeBxQ4rStcejaLdqNm+EF35dr1BChCYzruMK5t
WN9FbaLn9vCix11QiZ4XZrkwHppsyBJ5MoYgLAOWEkQt3BB6jBNT0N48pbCfFwlvhJYyC8MaACxG
sHxTV71uV2sXAVDgA+v5L7CCKTsSaV9dxnD8N0bD3A1TAWxEqW/tBTz5Va1m2DcgDpLaEFK5hMgL
BzjsBmEs9qKY5n9xjNPe7CCEMD8OZlKl+EHoN68WFZRdwkaCazMdvAcSSqbXzWT6eWhf25gbohG9
09wNP4h+TMP6yR5qC/ly3C2oJ55ouLxJUwiFXwWF7W/gXunfBFEXzOqBTnFtt94sYxl986wN7tdf
POSLXx0TrbwrNaCXZX1eBxeKya5gScxdmcZQgaLWjKYVnChvccoV4C+Ek2g3xfvj+r0xy0XPwjyA
FkfGjKZ59MG/NzZ6f4FiGkW2M+VdBmEgyAdnU5w1HtDOIFTiIUiCnPsCnE3DQm2OSPsfv2CU9v3f
4+Tr9/EIlrwsOyS8Bj1kvmxNVfQ8wKSa5AcWq9RiMG9kw0bOfDfOXksbeeZuyZmPDFpy8+A9e7LK
8t7IXfLoO02KavPVb/J/71GWFAbtLVYTSah4YF4ZbFEREPn9pxr5CqnJOgrKn5e1jh6X+Ip2ijXy
e2fBmNfRz0NU2W1PaBSHIc7PuWNIPAUy9TrJypw4ydb7fAETILY9TTPDhFFePTm1+Zv+eLd1v1Sq
DIYMuC559y6ffxE0VQoAAdF2XHvQ1bSfd3tDobYf8xM6j+8fDd0ZAUTQ62tPn32P7nQpLtb9Hz4n
8nxmEPoio3F4hPj7PZUvZhP1Ghlb76+YfEb5QHYSm2dq/pTBqdn4VwqofaS56l3PgGTjmh4pgfCh
kdDqCIADt5AcEOx/P/h98kG+jnGLh/NuVWobJYO4MsCiJkYYdxIrdSDLyddzMc+emqlWfNJ2hv9V
Rf6E6ismA2N5+v1oTXeclvzLchnThTCyAgnMTrywy277hkBkFgBFWuH2KveLXr96UYAJbup/giIm
aQdJX1UXL0gOAuTPPRsazWn3BoxDaIXDfuQS2UBlleB1sA6IZDLFYcSptVgQSShn52dPLt/89FBm
PKv2screiPWFuBgPCwiOPf99wbayKK1tWd+VzsFHSxOCH+mMw0KrZdEvDoC3pdE8Suln92mgQ5jL
uXbpOWANvV5LDygTl9aakQSwUZZOr90y9oL4MtkjW9LBQfq0upztWeGhvBAqZ8mwH4Qrg9TE5gIY
MrMJ4bUhIdgqBtAWBAyKPgy0t3WVbs+IBuI0sWYZ5LzcrJ1t2HqqGkVER/99rxRzO8MgNEZbz+T2
KTqKXyWPI+RK5dQe2tNIvnhSMFaF/m7ZeyMQyDHvjttorgRQCQkVOSKxn3osKAVUS1psRIX9H9KR
I87Itaq6rHbT2lJGOdpVAfxsrdYjHMUqGJq7EwJ6nkLxHsevHViIFYysCGwvng+JKnX7hlc8j+z1
zyjbRdVkg1qpZ+pkwGqU4vCYsB4emU3HJBJ5zuBBvEi6u9mJAELtrVjkSEn5oG7Mn9uuOgN3Ln0A
k+LqR0z5pqWDnePFEqDLL+KF3lOtHhJdIo5WB7CwRMBVcf73fqIWKtAYm8l51b1VsFP5dO3LpbaM
E/lXowrQH6fn98KKo/NRz97adlRzLmAuOBJUoRtLk6F0reKDwlruHyZ3SIbUzHxSqz2iGFUyXRDt
krLiQt3RRcelv4JjYGOJSJ9FcbvvlOUnulaJlQCS7XbCk3w0wlh1MtkDWOzeobBWZ8OFngEp3BRL
WhJToKPvDm9To+yvFAbksELf/Go5Awo+sxUpEiJ2qtm/y/WCeajL51acSVi5DqDPwbyRSVdMJFWD
Jl/OHU+qOdph3DN2v7Uzb8FvkbAiqLwDu3a9xojAm4X451BJXqXCQmornC88S1dvAZ0Yb0twahkZ
rEvKhayT5AQrfypLh6b1aB8wXZznqAMTLBS5LDJ5+PSQjIaqcTkyiLkruUCb8I8sLm/N8aRGQrAF
unTqC0JNR+oLQYxQ95VKtu9yrmp9hx+AjLjxiLP1pseAk2ZrleXMz+EaRA8Z+SCYKaVsAwKI55TU
xzZr94rwV8VpHgNo/9+ljkWqOnUTRYF3ULE9uEZgrvEp5dHsm6OdqApXezDsesRGEvDpocWSSt//
7NEhzyY6sNqNvSnolkKlMQ4m0kDsZnlHy+bvzLfqaCj5A8CDqijqbZC9htLEp/iWzEgdV4UJavuI
93sDVNHCBe2Irvgbxy0v0BW3PIdC3f6y4Q+r46M8q6t42E+QcsR8sgQu1ih9qcJKiek8LkH7Wuf1
Wsp6BggMKBcymxcGoSdVGN+fDXbg5YiZZUOha5mB8cfel6CvOQIBCLl8hAqrTdrad8FmrsmaiDQQ
S5TjB2TY5pZTQxuv6BoPU8iHWvdVfr2IekLkU3aAejhkpe6PjNlkTTQaT6JkpTv8QQgY5xzXZqP/
8OLRUCFZ6LBNM4PbmXZwPQwQ3hS5P5M2V463h2ez91+KjC/fdwXx4P2drTcZw/6AC0up9d3MLA4U
gBzbJVQXN9c1D3BPYN3PZKn6jjEc0RNWbJWs4gqo0E8MxGcedk0yP8RwRQ2vtaeG9iCiouZdtMTI
BANtKG0K+WkZunmaaWX88L/qijlVdpHJGY607pxbWb3wTo2ptl/Ml/XiYfVZxACdh/wDzNxSfK5P
RU86aSehGmWx+bhvjld34oeWlFPCf3rxoT/S4nTE1aPGLRgE9/Uol/VmtibU0uGcDU/3mXak3dTy
OYqv/bU/xs5u7Io6VcmjaYIcinmWUwlcEG0rL7Y/qZ6UAPHx36CL0UY24BaO5qoyeRlMFv+JRzsJ
fZLavQbj3SyhW9OxK998suPmeCj1MFzGnT+h5tm04Rnbk6U+DE0nzWKiUfDLjmiCFcTJXqu0o1bJ
MGh2A6M8vahHTV1var6OetIXQbf0KhtTFO/Kz3P+G9u7nmAyxxirTX6t6TI5EqmWhxUXYnR9umn1
ToJlGXXAYMBW/jZuDyck2+Kn/2iKmFnEFmHZPU8Q4EKXRTW94iBNWUvtH787p1nGI1fgaQYuosKx
YZ2daXt1f8VGdo8Z7ZZC+rw4vXOz6G+Gp44gYo2Jb6zk/xEV0PBvAgoHrnzp9iauS8ykGEqFBiBc
YbVB+xRGY3CevEOVdQK3Jx2IBRJF426KOL29T5ozNWxKmaiwLBiTrda3B6LeK62pJZKEWTpGbAyM
00KKpdQd1HhsDR71jd9qJcTZ5bckHaoZu3R/cWoz7kxe9UdWY2+xlO0nH/OEv8Udwtv44q5LODHQ
uUZIQ0D7+AQIq9KvDQnLKh/UgXRmngrjDTvxCVOq/T9rsfK2HyBeVeSlb/3owpQIuYKEdcRZ0moG
Vdo/1djqSL7cPe0NoUhCjyMSs/NJlknfrefG68PjGrWt+B9RYk1pIm+KmkT8EPKW50SPE4tlEPSP
n+HrcM+GMij5ekcWarjn7Shfkpb8b9hTRITehWSij2MAGPjec5Xdo8OGa4ou4lHOIp0lC3EnIGq1
FvIGeZcHgJxjTyx27332De/isFeM81DFc9fBjvCDkSrE7FnytCkbTDrvcI2O/71tCVrSPyHC3uYP
jaI3/WjjefGC7YeS3JU2wQ5HgQ+P/QcALpMozrACWRmbGL2lbD5Ha6HYiuqladhuOH8YYMMr07MR
RL9n9u4DGguleysbIs4S8rf6reQRR4qk33vn5IXT3LDGGxUgzit7c4GpSj14voSbC+ko2/scKCwD
z20BMzR/ujkgrbp7zMgWsIgPDpfVZavrIRdKMYGFqvArirbbapRbJMNi5LZu1ULfnRBKh13Z5J2d
Rw7Vf749dtyRx6/i3ZgM6oNFC6D5l7gdTL2Ym4LIVzOeAmJh7PhyjuR+K3uTuDbG3UyQDuGBnXId
W99b4U4Wc3Ek/SWEHBvBMbuth0/NCigen5rBMgHReeQsvw74dpWaNk22LjjMfM3tug239caTY760
Qi4YF+BEpTTFM7dCn7ermGHqdPmHoH6TAThltT8JHyG5zsdLmCSNMLfK9gt9KMX2bv3QwBNyfBAW
jYk5gXcEZAXrtAkHbEExEcO/CJZvoa+PCRcO8nzHHpMIx/AuHuiXrfdjSTqqwdwCvgIUyv/NV5So
2kLZGqoLRhl9Vk395JxRIsMBX+fpdaAw1GlDNUA0fQAfC1b5AgUrZISHsszosnaAW21fcE50MGXd
buzBmz/kTz/olUOsY9OEWt+aQEnL/U49IrYMSxMh9bBXR2CB7pifF55FLC21OiSXhlloNkahFwq/
yDe5CqXNy14ifeq8YUX4IuO2IN+zB95KXbnuIgzZgXN3TLQg7h4+aNBIbOAMUj2J5Kw2iOE5wGi7
fCy10Tz/g9r05Qe1JtzivfABGrBDGtTAFiINbInkKEWxMhdvyl7MP4BGT1rP1sQdtmbBbn6clWhq
J/w+Mrr5jSp54rS5Oz+tX9z4UizS+SsdkLutNRnQjWfeBY1lzkyLu/guzSEEtGVt3qFso6eqmkCY
Vo9tExmjAdO+33j7vk9/vj18YF0omzZNik14A762kRkZKNgxPV60VtEJ/MxRllp7gGU67UjRSLd8
8KH1g5Hou4FxK4Y3FoW0IyZDtfzqG3FLdDXtBUkXoyS+14i7Fc3rXpVSvwGbrjb2oXZquLn1msb7
TeYPTQjnTO/da9ZPW1e4eQFpsp7UIb/ssp+EF4efRKKbFR4rl6IdfqxheAfmn+Ps0TMuPJ0onsFM
TarPgvPSIE+yQaa5UBnXPQoPDjPRHh0GfK2yzqHzC2+h0GlGb6QcJ4lgICV3t8qScAnWTpVI2Q1I
vqnjrWTcAIibwdv4QKiee8GlfX1CkiyzIuGmAF2Q6eWwDpEnz5K6QvWUR7HOQkdGRuR/gb1eYlmR
3NjeglgX0R1BW1SDDyItrplp43j9YBogqM4jUoHppwRtI+osLFyQCvVSu+ys3i7WxIqgLZVqEh6O
hdOguIyEpfX0zWliu0SyrdifKaYOf/1ypMIA/79W2Ltr8NUIipPPplFcP7PecZvX+6dBCmm19L5g
a1Wf9J2R01fsOVTM5YxTEBqjAZtBcn9M5MHQxu7ADmy5urziWvlgGTh3vkUvQtCPO+EHsm43lQUh
/XeBzQ0C+rpDxeoojXV0JeyKUNuZ/5suwBNSXqTMZ/LZEio/LJm/iT8JNJ9gO9EeERcaoFriJLAx
dP8AB/km0Bp7/xD36HYYVBWyAH1Nw2wt2amyUsWBt67a0ZQNkrLBtnqsYm3xNJQzTJWH++IzeYAJ
EkrA657uja4SRJYHlpckC+l5USl9ZfI6wjJAAGlWKFBHQwruf0Ad6ktQVpM2gnJ4ob5d1cFUFby5
pAUoDMUcYoVhU0/Jkn6S4XMa1HCITq/FTpf4flI/+4szPReFKqIcRWeUL1QO9BMFFVjhsH5QMZdS
Ia08kZwWc0QHizsbDuYJMfs1URI2mwOUPJKe05vxed7fRq+vzdixrSh9GrYtaGBwKZZ241NOQOCF
7NG19vZa5yYmDZTR+Rb5oB+HniHrW40KYPCPqMHlqw1yfgQxcmItUf81MxMulrCDXzbqn36i4oUN
lXai/8OQMM1iKNE2GsIV/ufArWOUgNuV2IlsMGynPzsy9z1oBaeLMZ2NHyPw9Ft0HQhvy4R+K0ay
JnrW411gM+XgwSGVKsAcrpYaldfuYtsYBSaDfrDzMlPD5o5KIzJmrlWn4bID29WR0wa8yp9VSRWO
jGN29e26XmOxDfe3bWrMONgpWIKVwPagnszVrPvEZoxYI0uPTpZ28O4+24HeGim2cAoSixoeDZ28
+wcBxFOO1ArqcIgs+Yf57xYRGUNV2ISIRylEsMzoSUFjGTBaTP+4iduGHOncN8ARwVv8mX0sf/R1
s1H7Hl4q5XEphpoRKdV4+3yTGYBDEce3ILPDpYFfeFIGaa6Te27MYPKTf8ksiO9m8UMZuSvA9H3/
dKRqPcZVtLHNk73adTdSnUYxfi0TlVLdcVPIBXHxjeIrA8JX/XGDDwxv8BwWMNL2QGulLiCF4fXF
7Dzoz+WfHDlGhSRxDOGYgxQxCGHxOXtsY4XWLZphpLjS8citoQJh14l7WM7BV+bpfbihJp7Ompqp
+8wPdb7bL2QH66UKz87inSg1kVEkFt9RIlfdHtU7NeG38fZjn/O5KdyP4LPtUSLtT5BeN2kfSMlh
uIga2e5Eu0e/t75MJ4sSDRJoixRfEHoQqjIMRjMD3CRiRKu+XjtpIJ51bMCUuICr/sOByPZJMD6R
lSX408MG/pgsdr8sclqN06xU69V7sa8Zt46up7Eg6clQG1ByfohS20MSE7iyKwZv/i0mIvPWzVwN
AbJnBZRFfUbw87lgVvZjQE+00MF6YskHy61YF7qW7VMkTDo3kpxZT/JHsMg+Sv1jXl9wDuHbkLKZ
t5WBa2TMrodC6Cg+kegq87SePyyxS93IRvsSlcdTS4vbQPIcWcAjwE2U5kPb6qY1EFyaT4Wja4N5
LQItY3HExSYgHnIC8b0DL9zt0W2S/cwJ6FrvxWBebDafEb+dlxHtmtXx6B+qBFzgKi/EMcnwMdMu
1cURTj+NTJPTqIgrl1VABRUW3UFdU5MN2DwWdA8oq35uFol/iKdAM51Ny2CTAO0BwFMQCArODBvz
+i+W0Z4A1X6FUGAN7kpMM5P8pzqznk5Y4u7vUHyr7E7+FWcpCpMysFDwVx6PKAHj/0q4MCfX8Tw3
8PbdcmSL+uk9BVuEz3TfGgd7fh4hIP2Timdeq61cLGLKLr7v5K3oMwGX9FCdQNhsEjQP+pnosXQ3
fpJoyxM7WsbzQBXrinZfGe/lx/uZQJqCTjMJoD0NcGffhx6wDdOXKzIMGMnR7+oYVnL3/FFDF+ET
19UcLcjpclMoZeNha4H3LSJI2abtFBUPhCeNWa+G5i8+Fjchp5gAxfXrcwpBUxwC19GE2EK8J/qH
Y2tJ01vY/XMj4k+XDql73rptwJpNmC5lYXzo4sA/xhr1DD/ZWGKZ5zlVRA3GMz0jhFq0hfD8qI3w
mfXfIofrOJt+ar4oWxDOBghpXMRTHTVFiDh6oA3n+NQttv1N1nhd3Y4beSfp+lTKA0ngkPAeGJDP
xSBLKAwZrCtFHBZYQFp60/4uPobW9p1qTN8y69WIAGEdCGcrAvPdI5EplZqBSfsW0BUDQqmgTcpY
yuJUukctD1Vc+KYf8yQ/hFkZmlC7GFSrt/zGe/WHFk0nn0A2f7A/tPO5Peh6K6AQ4qZ3q59mHFVB
C5Z7O8Q3fkR6ivHzv5Kdf6y+UKaO4aYUeJqhpmZAv+E05zD76dhltNF8dbhz1hcYzI6F/Ju1htFH
BL9/rDqEf5DToqtTsR1q1hGFi2Ei6ZAPnfZL+aMY/jdBpaCGvxnD6HWE6Ls1rKBoaVXc5G7Caufj
pF1komsFAjkqzYa2tJQAmgUgP0/Eq0JwjbystJljGrTyCEgf6tL2+AI6B9+EGny+bFXGaq9pZ9S9
PRfOhnSY5L+LjyGmWKy7Ve1D31Jg93OtMsWwrMk/jB844SHWnBhBS/ZEibckaHIjAfcIRVi1CJUo
3FyO6UyWxvk4LH6mDDdpokB0TN+j1GCbWQwtCpZ/kmdl7PgR1yLFOWvFAuj0qLj/exBeuKgxsC0i
xatDpAAugFJ6klaLQ5Dxq4uiht6CYBuZAcXWnuY58S9RlPMFiiVXyt+P6xaOfVdsTWbZbcrbISKO
z9ifzrfnL1miqCHbwo17Rx21jP8wFl29boetP0BrlqsF4ctRsAoeB+O6wSrwInLSBWmBarlmHrPo
z5rMz0Lz2sPr8gAZXSgB7PGG5TXB7m+qfikTaWf2RtalJjJbDkeOiQfCeBGyK+I3A1ywZwbTTURj
lHZGGObeGTuRt3dwxJZYqd1d5xanuBEwy3Dp5UtFSO1K4j3OjwpR77sBKjqTnZWYNt1obGpSn3Kh
9OEUP6HvYL7ROYL8NOr/XULyr8Q5tylZA7XLQi6DRnPr/6x73Os5kOAsovSrtzwruBvMh5C+P9ws
e+HRz87CcGqcbIZCJsPYZlAl3xJWN7Ep9RLVmUJ3Lf1dESKUNI8IehQ9xYHEI8sWkzRkzA4SjG+E
vwSrvpX2uYhgl91rkFyqCTj5A0uWnJYeZTQ+q2ttU0lVSZmAxEYm1dWkG26aCL4I++fNoWDA85Q6
S2gnnkLKeeWKye4ylZdwplh4MJ+G/7R0n5a6TOPSJeDiwDdrd6jy4LBAMmTOLKy3NxTiG/ue7HMf
FhPCOKghfjo8WnAMcEyxJwn2UlXuMvIUZMTd5/oylmTexYvsk1HjfoMU2hHkUztbgdJ5RpwWU3cU
9ANrttvTqJQrlSK79ctA1Z/h00JpzOAqTA0oA6mfG9jM/iShpysWcpNGy1K4PiuHwlLXeVNzmmQd
5nR4ltlHyf9t7pbVXwWwudwb8wjIPe+h1mctP816KEqd7Q6OwIrEHPwoOUdxq1OypOEi7kZcV2tV
XaYCmtPwKPhPaWSrikhknuMFLK2G7gRgKvlcqMw4Vp1MUp1lrjtfglx0b9+fF8h8RN/GxK0bmsjP
rtAV3ZkqK0/uR+jNSXpbTJ939RoKy+QIGLvo4UyWiVF+EX1tBHoCIdWPGgALECxvGHyHQjOdDyov
rTGaf+ApsXoVke0neD8TiP0ZcvZGvPfXmW1A4DQrC9a7EWPDIMtsPBBwhKdKZw3BJcpe5Me59i3i
9yV7N6uFebaRjDWvSQe4IAWHAd1wvq7gHlkYFIQh+bYt+jkImPJ8TnvUb8IMm4aBQZYF8oHFH37X
b+FeHuRRAposm3BxbQLRQpBVyc5FgAhXGz0nsQq5bhBWiSUaFHoTMyFgZO52R4FPpFKbs9wVAB2F
hUU/6Kk3W4E95apENgR84UaGoYmqjsJp4yuD4LVw2Z/Nt0FoOzp3QpfFl8LrYWOjmSbcTmk5eiJB
ftowkjfpXsVmDfrhcEFvrtHyFBppAEf3fzk/tBHyEOIJrLbi9twp5BOuDo0SOUe0ksch4+oMakAL
xz3IcvxmXDxwu0bT7LaAKt1WUlUH0MBaohgn0l4lRvoRyUIEoPrNiqBwdMJepeoTXNTFNcHQCMnZ
yFR6WUHBuWHj3f/IiSm6ov1TZrB6vwzT8zX8ZdLB4wH8JlOiH9x4fwoqV3nV0IlT+nNiz8yZQq4y
nFixGeb4hvuXrKIDxJ8EyEgzO4pNJIbc/qQMOFjs6Ir3pS8R7iJgyzjF/TlX1tYc2x/wL52T02Ol
6+K+g9mdaa3jrY+/UMteXf2T+9kIxIewp+yEywwMX7/wPw8UvawmJoZx4gJpC/cr0DdAxOIXDTPz
N+Pdx0CzUf/FHX0XLENHe8ixIfx2ATNPYb1Afczt0MgLxZ9xx18K3qRsJY0fxqe98XG1BdXzOxVM
uQCguPZQ67I+7L2hYXCL8+QfPNg6rQtm3nsL94xNrCUwzD3a4kgf9TAIWAJZ7T5jLQ9JOIEKI9hZ
R/ZSjLmBiDQ0FRnzCAeA56HZDuQA3LYIsX3Is9PSG6JwZup83gSEvW8gvaWY0T0fgfU2cSFY+WdS
8UlX2AoonmiVZulaFJIcwzZ4xD7bRcdjJZIzUKA2aASc7bnxtBoigFDkkutaU4eAqxUth3NPE5Ka
AIv09m2bsxw620z+Hs3DnB5PrF6pQM8sDiNkdf0mRRG5jb5jzrpKd7p6qAQ0pcAoWynOp7Y5falh
gO9lUEMCNimmyb4z0bYtui6ejpE5P9FP2xdEDvmgLrLGswZs+HHwrsvwOjFpU521yRAL7J/7QGO2
pBmFmnLB5SQrBtk6vLnT8j8NxE1PDO3DLoTtjpTA2oXL0nDwoVHzivRLJCH9zlVMIDpgWyHxl4Mj
ozOBEaDMdsR2HKC7YgDHwvc4la8owCmFkw9dMnvMlnyAA8J+0oJlxet5T45Bg1CDvV5CMvJxMrp6
sb+cspZJ1oMvLBP8Yphj7vDMD6NFSxplqXjLMEi0odh7oLjMovVaomfjAtw2szJ6yOuR6sMsWyaQ
FEqOK6FbLNNJ3dPnpmLSP4vllt3Y2808Av0KOucKhxzR3E6yJVxH5OiYVruAtxxwZaGq7T4vjdW8
n8Yy7Xlw8udvlVDE07O6Pz6ZlQ4n76PK2x6+jwv44+yO55GOEShJXNcju/prlYqJgqfjHjGDVolP
x3yeHMDs8HFU5xKBmW+PXznj0yjne0taB3VkwW7lFXG9h/6WdAzBqxiLdd0CCYUeE643E1xG4sev
gHjyjrtIcNtnMKoNDDX5GULHqOv61lfHV+CU07lXYhxIYzTHrhp7ZQ6PnW1YgE4k7wkYY6zkmETq
w0ufAsjcEKZkZfR8qvFlW3jfkq3O2wPqMrEuVrQNcv3tTOypW5oZnEXK+c/phgNAP2p5KYbRCLNf
J7Ya6Md9jG0YZNU4Ot/2qVJcnGIBlwzQx2X99LnmV5ZR5u/KMx9bYaIw4jhnCtpYGqv/XQJqDAwt
YWq2WKXYhx/M7bHQtyq18AGBVpiIZzgWPpXQ29nXIiW9q8/LAssnrZPoksXCtMDNJ/q4OhC3vBcw
zQf7hFm/em0DVXZFNqu1jzwYLNZOTx/nRKf761xYrZKoexskwzo/+2hBqVXnWS2jGwIAT4M9pqtw
csZF/1eOz/AVXhuDzLW/HR2Fzu9i2+1BOny3V5LrS4syoykRCErXXuC9as55hHmPk4OzfD2aGN/+
ltWRkrtSOKKOd4ZSfd+t8iB0KFYkGPh87MZzuTNzSV5FxZA+oPRCvOx9w7CdFD+BkGd3Z5DtBXhO
imKEbyC9UoD8rSDdpYAaYOC+TwnjI6d+mqzWm62r58GQb750ETks8mc6NIYK9+qW7J4EUh5K/6i9
2S9zYgZMZYig3/IHyBZGeCQHEztuvbe+i3t26zEpA3A/Squ6h7qAo3eIEReEteqm4GNjBhVaWMEn
jQHG8YxTewTVuVANdhvwpw70PwPAlaP28UWuK1+YCvQSO77D/tI7Bkjkry6x9d4I7BN6ewAHZQ4+
BhgS5QBwDs1PVZ6OILlHeiV24JfUSljVgo1hnMnuvdhxxLPgtv/XKyYi9q7Tj/k25EEwW99c3T4E
jVJvgSODUOMmzUEmCcQlhGAUUfOqjA9tevTzVA4umK+OmRqaulYfNoIhNHBQYt+d3aX/6uJBBn9j
YDOp0yBACDdlTxT10+kvgDMDLtCBZweyv0Rzl3wa77Vq6N+FBAtyNGNMbeudgT4IVe1WbRbOPHl8
vOuvBdecJxaqiA0eaf7jvDO+uC1qccqVh02aVmCK+IQAi8q+m0D0qvoXS9J+vALSqdOrvFR46MSE
54wi4GPWVdVSW0MJHxbdQS9S43EPgvVveCwL5z85PBrgpZfuI0BUx19R2dshtDNOOF11aKfEhwz1
4sEslfl9Lam+KZbyRpq5m7MD7X3jknCWoSgEv7sclmNn7yzeV/VBe7b+ypUtQlhhWknFW8eJyWDn
pb7YkgjCYNT+ztnBxtk94p24/YCm6FAxZ330fOJyXA+i8lFPFzynlW5XoLZrAYQ6Od58wxDep9Dy
k5Jc9tQXpRwQRSzDE/UWL/eVI+ZIrRhlnWpxWk+mYlWNsaupKQuQ9jcC9tNz4gMRuVfvAm7131qb
boj3nAJotwuRbQ3mkAdbYKaXWK6ITxw7dUpGRwRJd3euEP3m4rhnKsa7W0njYqR0EFzWxVc/m3i+
Xmwi3XwQOD62EmY2jQScE8VxCSCLOxPQnLEFk1QwjYjOjQi34ky4CWKh6iTb3ijKXcEAptrB+FPT
GAL3AcA5JK2TWTWoYTlqL/juqsGhgzLK4xPxpfdTn0qMB9yJi2uaaFxF/cYKWh8ktd66NrNPNn1g
iDRf5+Qhy2RwaOSDsi4wPekJuaZBQJ5br5Z60Mt3HYLbLjPkswz85YiA73JYiwyqoRV/cMiYtvKW
5H5ekeKZ7tr/RtufT0AX1FIWpklOF0rtMASQBJCaIlWF40aN61w6n00Fabqs9jrvRVJWTSHjGMQR
KphWILqk9AcQuDc9HYGS18Hekg86h998VIQrzOWEsssj91SFoQGJt196pzSFNyy9zofvfr44TpkM
o0xdL16WnjVDA+kqycIv9+hVmJ7d+PhVbRoU9JHBLI4UaV2yUXVg2Xh89zARHgOs6UeNNmMCogCw
HFGGF45dBWt8H7PNjobNZ6H/fuL/WRZQ9rxUaZtsbHZ2ODgKd6jG2PupQ71welZji1BvSnfqyTfB
9eUvzOFJqUcG3469LEHQKZVxZFSu5xvdkdG1ViYC2SlG3wVbO1rqOtiE8FM2dgnTp8F9i9fjpYVo
5WzxTSQorGMTDmmde6ePCu7V2x5tvf/OFwZURcleb69nEq9jk+GCCtK2zQvlJAmKpaffZhHULsdy
BU+xBgcve7oeUJs+hkkDEZLv783yMNeAyaf8MpsWmAfmyY15iT2RkhKLOe1b1M/3E8fagsjuAmrw
LNIMv9hIHTqTdteJEIo6o6TuSx2xYAgAsizq5ttHo1FtWwvSAt93BLgk+UciPU8DnGevZvgB5Wwm
Y2dldPuNgkPMrHnbYi1SDx0ZQZRcR6VrhWi4WykeC6uOu0Ti9ooEXo02d+CP8Ps02pnqmpoL04fJ
vSSOk/8uNo9h/WG4zSGvx0lj154yXE+XoBa/P6F+HWoGC4We4ftFIr8ePillfqo/pBTmv4uXhjIa
XOKW3lOTCG0LBmrHZqlvHs6I0xpkXK9p5rndqpWLZ0BELJmjjvi1filRgzdgIsGiBhyTUotklD2Q
OkRRPPo1r6SwSeVLWTnOwY0jbYWbtfR3tb39I3TQI/MWBou/6Ump083srGQ9V0Ci8bge/y9WDm+u
EVJAFe+eeHZ4sa70I3qRoPG9x5bgR/9A/9n5g1gV0RgTG8ULFdtdBVW4AyM5XFmElCPnYkhKxngj
Rc6tu7QaLpkjpQKBJOaAcQqSCTVOpbnjv2jY+Yndb4gIOV2NqTiklHjVHIrSAaHPDmJanJGbxz+y
/V10I9zQUK8lyFU9m7RYlK6IIyxNuYx5wuZa9UuFQMAMlXeir3cDg29KD/+eHP74SUj0vaFl+t5y
xLkdio996BBEpGCs73SSurBdhPpB5lfIsu6d5S5+iwdR8iXF3TVkyWYa0liUYyOUR+pgz/x732CN
6LFmQ1p/MICwdXQNXlwX4JkZ/hOlDjtjPTOAgS7CwLZXTDCkiZ+Xv78WxF0Ct/bHbfCSTDffWkA6
sG20FqX4ltC81EvMDAewLWTSMklT80Gn1S0OGnjZTCAMMWjoMUxwDwAmOVU+tJcZllnmsEhdL7jM
WbJjlqunalWLIg1h2zWzz61zVKbI3NSK8eFQQDLGI9eKsWHH7itNRXSz2LKeFOsqNrXLGVdbpkuX
UAwzolMbH/nuNTvvTRjzsn5xt2o/dZ/kl3S1U+VEplSAuZYvne9y9bLWL0Zzh4MTufBlFjUxz3fH
Q5SnVdUgdsRMIDuTRSBZM+A5BaH35prOsY/dnyDm9TcBQC1iLU2Wns0JLE+aG+CInhcfd1naE6hu
e1es8QRw5VKd+LTGBP/4rr8O3wYTMwBucPPZ7h99TR0Mv7E5QwiYJ7IhNNu7XQrEOGHJWoTOKV1b
DyazWltoalxO+UeqTvjj01IJlkWzW40g6GzWQDW1VVBtBQ0M99uxdv3OjLTdFHNdnsngT9YB1ZEY
IavlUmUyKLf5cS2UDKx2EyHrdtXHv239kM/C8AHfwQFnTPqXXFYz+XVr8Tm9/xCPBDhUQ8iZoZNt
S9WN8BT7FdlluQoNUA388JbBxhe/KBSeI4MYpY7IvOFVP2KXZw6LP8Kmncke+QhGCwpiC/SB0qR7
WJmcq/OUDbq05ICkG9zENoPxHkvbepTz77xBgeIF183Jezzb8lmwqiIWp9L58cmXqf/tuO37i6Mp
qZYqA4c5QBhAk1/tLZoV66REj1jVOFgvqcc1rk629SIE7MYHjRjEJHK/OESPRD2R310JCRWK7c6Q
qoCxeNZcZnWt09X/fcJIRBTE9D1xcMFFqEM5ayISW0ud2yP/DQO0px+k/5TtvsshycjId/qmENV5
unC3U92wDrRzlXrH2+cIBuMQtqS4kgUpE5LfOhiJcFz+gC3IZJUg3hFkezswT7jVOz0zduEaoTeG
EA3htLforrot1YZNCKDTBfoz8ZZXYGLb8DCq9reQhrsJMJFwW6uJoRiFgbf6N0Dae2cdgmStRX/D
IC+Wp9+buGdYcliF7vzxR4rNDM53FLPUzQohEil2euxe3yL5Z98IWGwuGlVl4cwoS90yIQeiPXRe
JbOywVm+YOkkfR7f2VRqNvCTkkmDiOWrE5jGxCdvd9yHSPRPXpSZXbjwtiY12pHA2+fJrtJ6zM0p
0EL94XbLQ65eJnbirAD8+pVndufbFrqj//fRUDYn+o09Be8caZPYI9+qD4Z9gZc+rDnjpyAZyXTs
GI02kEUUmwv7e1lgSmZNCIdjp9y6ORTXmfiOErpNuX6STX7QsB7qzKIWH13U8Y6abq0xDyuFDfx8
D5U3ZVjh03P9dKUGVTLg1YzTcX4lp//GlguYwA1Unz679U8Y+YsYgLkV6o2eYpa9cOS/uyYt0hHF
gK2VxEsTJU6NFl5sAL0s0wRoJ1nF38r+NPUG74jSEm15p9YdoLmc8QXGV1KDzPqqp6TYMQoRGk11
6tH6BHCnLKASvoIyWHkCW+SQ73ZtPm5afCQeUEJkIYU15cMb/5+RaQR/+ktxOqPbJjPZM+XYU9wf
3Z2h1tRFdSOUlzswzZ+Q/9rOdSUIAs7sEtsfIwKYbZrqdnQEb907KaSeI2ez825ObP9RJtL5kl+a
HeGHfodKhb0/ytL2icPbOqNQjwZQijhpAkRbvtQdNbO8FoyE40vAo+6n92G6jnsZAqLvTIah22Rf
9qtjYfygi30JNWt32V1uZDZsM07ZNNh/l/EA6j3F5LBXQlA0A12SdyU7o5MYCF7fBJ5YsK+oNm10
BMM4bdL0Lyke4tZlb1L3lPmbeTnengOPIboQbelDEAAKeB2uLJyhF9kWrzdCwwgwcyb0QXnzBEYN
++BKQfi6cjeiGmbnVh7BtncmiewAHdiua96avFhgH5auYo60kxi4/4+vTamadr4CeUAiu9szTp/v
ls6erc/CpI4ziRX8OBLSsD3jPi7VWU6k3xrGRyFkoeMdL6lkCqyEitNaGQzH6ketXi6x0WQ82l5C
Km1XBluuhlhXqbUkbJm5sMpgML74s7wBwOTcjhHQGeUieDRI/fLTm2NC6nvaB87nfXLJcXhbXBo1
ZO5/D+1DlcRjfLzS/Vox/Vs1dJuFXnYU2eIQO1xPlUpBlzsFV0U4OqfJaaUc4bkz3wiZnMn25I32
H1c4NEgNIekE3ix9iMOCuoZKmHlz1wa5lvhBsoCLkpkqX8+YoyPqW6iyUhBU5rGygSSZ47vqtaGL
HXKcfaInnwNynPQb4bxuVFIBGTwwydNaSjFqFzDQUukwbyG3ivhPiH6W3Mcm9kPcuzdtjxDCm0vd
W1DDEz6+44Rn2f6k4VDdIQtkdSFXp55jCwE82iFI/LOWL3GwUAlNJ6rmmbjKQsOy1zBn5Rw1Zyux
XcOmdFX9kqMwiAWQpowt0gxa3l9NNHfOVwd1UL3LvpSa3D0OtqMMw9wEjLG0jrjJjlfkrweKizn8
dhyhGm7QaYiGzcbwwnsnKQ79OtbO8CxXs9HuKzfiXwc7Ag4MYIhjp8H2rooUSRc7dlQ5I0LsJR1o
/VQNplvXOjhHhbGMaguJ7szxIdOikRlAiVzy6zOpgqdjB0+G/EUPwDpGc0HV1cv+OZ/gdOgCYpb8
RY1BUzsRPb8E/+Q0dAEhMf/x42OewEG/WypExh8braAQjLnEsB/omRaUF6EW5ME29ZS/odzkrphK
TpZp3s8F9SupemlynAsdbd/MHJhLwaFWERLW7522xzDRifzBnc6EKoqWLpdKoL/n+UALwpg4WslG
J6wKTxqQHoJw7a4mi7on9TJHtbbHuAL58dIxVgI+7EvhSthwM+b3BSLN2/Cc7ArzSNpAjooxYkqu
TNnAxIwjHCJNfJt4d9+wZ2md4VmGUdGV2YadPArZzCRdRrjjA936788oqx5eD3IoemwPJkObcGBT
e6Oa8u0Mr86KjddXE1mFMX3eFlm18eyHK74y1KalxJMQoiE39g6URoS3GKVYNdm62L2NEsS7v5LK
N2/TP+hNBlXGv1+a4rWb6F68iB9zHLMRQ24v5KtChRBhQr9EwDIO3i6MJdzeQDvL8xiGwtpc6C/p
pMuqKp/qj0E+DN+tinRgRjdSsBU1JBxh1GAOpD2Z/NVQKvEMKFjbYeU2QJ6yctHj7XfaNcTINJb5
Ccjmus56rDm/gpRznoXtoFFAbN4n7zIUeEVJ9fUltXjFw/kFgQgblLadVRa1kX4MsCwn6+mlXeAT
+ernFq3tRdYqnZ9mNoRGTxqSKUnhhp/yi8IBHyPp8SJkNnA2P4ve8SFQr/XYvBp9HfbZDP6rRLaV
TYvf9xxLbrzV9UHS2zLhZbAj3YgY9yyr5csnM32JwfviA9tszbuPG48JozhfpRWFHL7cf1ODbVrC
QKA/AyMEJO6YmGrhPDxPEC1n0hxZZYjy7jfQ1vQV1YfxV7btOOr7AamDP7Wk+RoAnsHcndg40Tzg
KTnoBZKwNXUZx3iIrc0dxhCqCKUZdM264TCXhMcI8mbPFdbQ7gaSHFilYO0qfEtFz76b4ZyKXpt7
5zAZuleFr+YsgOl0Ud8gFUjT2yB3b6q9M7r/atDF+hknWBfCzz/bI9DWWnMfudMF3lqQI7JtEpjd
gWPalpH27tCnm943zqxE7XTY/ynNeuuXairAOThE+6qvzrT6oT0MpN5fuWfBCgnl1PXr6jqarbnR
eEo2B2k1gluEJT/aN6VeH1aC9UoV7Gr4H1YipQR32/3Ls5x9aYFYb6WZUZyh4NhxgcwPPco7vf1x
Jv/xAPJjsJeTx3LhtyyoTYajY2b1JQRKoaxGe8yo8CE3K++SMhXSDMy8jIxcn3Wd07Tgq+6LWmrY
vxAUi/H37TwkkGUuUQjvJka4E3uYLk4XxTY9E9NEI70VpyihVOVcxYEIjVejmAVZ78KJDQHu1z/6
d+Xcj+EYgAQ58lX4MDV38RK89SgBIh7zXx2818MtsHX/zC1kGcMPhujZeDEcVAAWh0/d/wlHxYt+
a400UIRYGDSU5MwuBqkwavMziK8/LRwqNOhUxEpGl1SV6QozbqzsDCMxswhD+Ksi2iEx61kECyS7
IzAJ5so+e4doAlRdF11bIb4sw3F8X/+xvA3XXxRFcukGPceg2k+t+ek6B75YuiQeAl6QPWsdvklw
jH06j31KHNCRX6wKyOg7kLiY9ujhcvSCJqvndkwInx9LC2TKDUTQx8YR5Yj2Tyeld1agN5z+Tms9
e3yapDusGvIEmObD7Pe4ePf6TJHItcEQI1pb8MhWJDtJr9elJs+9qMgV1jr9m+eTYXyd88ORZu/n
nUAI4G08vWVIu2tpbiUzwBXnKQ2GxlcAeyNl+tJv/Nt23KYtX2OTqS3oi+oFBRAro7kKFQ+YaxM1
FSksA/622Jf31zb4AQqu+1VstPAyMHsFGk5rulNgeonjMOMKx0loBVrxPMlMF/ft0S+YRrkMnzBW
UK12l28zM9a+iOVIzD7WN+fOcPHSunxzeKrrtSAkJuSx3jrBShScbkwlDZU3eninkzt36qiPvohI
yDiJz+6FVzBKZuTAxUSyqyt00h14q02wk+dT54RYjC1yGf3wvWj4VG4dcQSkGkECPIfs7roYEGFH
l0pMG9h4MX/NEn0Ee3mn5szTzsZyLcOH8QRLRkdthryC2EuzW7nAJQDPpU077BLC7uffAEjeWL3B
s4Md6IDFhx4xjqHImqSJq6KSdlw/kl8Me6nnI9j+QWLPA50FAfz3/zbi5vYDgnpXBIJbOUf+DIYh
p/ftS98D0T3/nCCx2NQkRJg9mFYgbw37u8Jre8HTlQv/JFssJVESWr2ZRUc3fIqpQNDUGF3fXlZU
qLrphn8vORkhHP6gO7bQTj724wbY4Efu2rtdgWYkkHxrholpp4ew9NvynXWEKV47vSNUMoLX8vpp
CD50adwaDdAvQxpct4DA0qD5ZNmDUlaVjdzwiiuau47/E31R3gPMvP0HKvfShRlBYOq7sx6bq4Od
UhyQAPw1HOR1JDVnn34J0YbMU/DZxjK4mPCTByNsDuj3nEeGTbBQtJsAGr5kbm8O4AG11Q8/1F0w
OiG8exNQqhBh0Q6mnFIDqLZJqeoKquCR3Ek3VZVN8A7k/9w5Ljd84zmiJ0zN2ABarFQX+0pIBpd7
2BGyJq7BuHDU6gv7/neOAd3Nz9wRM+jCmoPpjho0Q7ROe9t3FAkpoksJA+7gFDPJHASenGBfCgYB
XY2jnEyPNafqAKt+A1VHxV7MC1QVI2JgJuhNIzLWR0iiYo/TmOpwY3Ndr51qN4qV2eOVT9PmAI1d
EzIIv27rAIuL07xfGFqOkFRUYRFXl24wLf9cRED2583k2BsHGPRMe2Wg6yfQERTZKVZr2velF6kv
80B7kO6I5b5L2Qx7JC+T4GC0kZw7Ky+scAaakSeTnx1RzXcxidvKTkjHx+ZCZ5m3RrsuVwxuNNPK
BGLtMCOC7uinphLTtzUo8rrd08wEsk+nuGQwRhpI2Zc5ogNNcld2S24hNVpAoV9QRTjAeeyt7lmu
cjaPzGwHmIwjHurAe6IySmkOoXbksZ63YN5QZZGTYLqwJWOKy10wteU+tmetXR/Nog5W0vuApE2v
YNOWr4/bRpUvPksLRtmm2uDctQGLyHB5bpZnev+YzYpQvq1hINVY8kMmVMWmjCpqJFt7WYA++AUS
r9SU1PjZIDwIbhx/s6zqwhd5htXddU1KpqMgR8Zxjv6Xg1DgOazSl7oC1u/fnsyictFhFeb9BPww
yNLpAYKIwSNxihwCNGieY/E4KJFqDHzBq14/wYCbOPuGOO1dCRaiUsgSUMC2HsIN1ZFqXh8ksfNr
r+ul+2CMoFHI/aRDgIcOt6A8KATjf4pFIuAOZVyGsNzOI+CSzE6gWLyKcvF1JjJTuMzZ+dKg8kpg
kjDo9b4xbydqhE4N1YfmE05I3I8A9aSwVFvx8ty5GeqJkZ0LhJHuPYEfllG55U2I8RflrVEqDlow
/hhmkqQOf77C8zxWpc+3xA1u7xE9Yt7QHIZdqcRToESjRtXM58JMYluumnuESpdzIauzrGmyGV3y
NWKBNTpHM2VYgIcz2qQbgtxy2B7tJNJw1tT/9vBMX2oMZZCEhrle+hlxz9eBUGZF40O40ZJu0Itk
V6BUUyu/nEqDx/NXqRBYzxD9ygdWxMMe7wsLcsBjc6coUg+YIwJOt6B79DShkXX8N4scwJUIAZzS
OLrD3p2nuc/Uv/ciPhq/yRLkeldJoyJKwIhp0QJUBW+jhkRoVWXIWHbHsF5JY+HBFMu2Z8sn/ubu
tnj1gZUAftaPWm1XaFbRysDJCq8XjFW1iIDAPZudXFQUelUvlb3XBX5oGU0kaO9RtbLwGJrSm2rC
3kfuROwzvn+tf4HUvKKdgIqoNoDQDVt17yB8/PSkxf6wlMXYBLLF6/uydp5QfKYXGmZTKslpfL/t
6eCcCaoDU13mPAdUWiXUA5544JEl6dxXau/D9SWPsqb21He8gDaCPnhrsvb+vAlGv/gmbl2YZxFs
kosQCodpotLzMKJdlw80opRUpPK9L2EL6p4Y1tgfUBOSh9mLUAbGB9/zPpwqzuFpHZLsM89lH6BO
VbbyiiyBLUlAExX0X4SxUgRAo5mdLi7D0ryw3e+Qz63R0munzopfDsAcLHsoGJevte5sqZPoaHQW
Lszl4lSlcHVP9HYQ66Kj6lvI2T0N840rTaEzZvYP77qqdsq3GhZOlIeb51laQ8gs13Amvih9oQG3
VssE5i1fYB1Zs+HpbGGsJMzDg7xX+kVel7huLIspRDNtS8uoAUNmZsjDMsows7D5h6QB5KB0YgxA
nH8wMvFJxjF8biGr4FCWDSgyr7XIlcoWXlZnnWJkk5nx+iHiDLBYxnQ6E5I31Mm3pb1NODgt9bhO
Ud9oV7jJE2paWiK2xEtljBGz7In0DL9KXixXtciTOrf5oLw1JtkRkJ0WBuFOv2hnTfZDPgGb+EIQ
emjJFDVoIi09nlHt1L1qYFEk09S0/EFeCCN7JziP86prtoyp+IA2tRCqKZdc1q0QaWPdbvdGmG61
VkOAmmN/mcL7X4Nnhas5QsOQBygCisvVBNYuYvpEwtFHldHWLuVYKEIpKY5uxnRkD+sA9avwq+S8
adSCz8Zkq/WuwZqWEqMYf/N2hgww58YyzvOR+oKjmGEr6w8pQiacpOLySm1xofs7BR5ncI5j91jM
2Wav6crtULJXIQxwThAOf2yZefOMjK9RlRbyx2DU9eB4ISnE9GUt14J4dDTu0QH02x0Jqtxo4QY3
jYXoVvs9mTPFhQP3dbkwVxJasRhdLB0Ch6BCJjkRd7BUpyR7dNYWSLEEXTdiDURtotGLINKNeU6a
7/Gp5S2UKd4JpA2XBgqaIhbC3AVSeSDVz6SlvPvJcvCdN2WDC0/TZlD+PYl/PLlh6ypAy6wnAUT0
oJm7mpBmDsUSWq+E/lyzsogjslLBrBpC8ED5KAgJNCaDgHITs2tDCH4U35QzEIdHvTW4BuhJZOWI
zp7mphuXMfvG7uVc3nHecd9BElHn66F34Ombru+yp0X2RLvp/CHzVPp9iuT5RSb7V2CczUbjpqNY
sT9CIEIYuGgDdTFawyjbaJqzb8R4PUQC6ynYmgpddsDL5mx/+DX/IA5xmqnMOHlF6fTMUFanqfqD
VrEpWcHzmqNiRZyv0BuxjLIGkJ94ieBt5gE9oN3Rgtax6uBo4e5iWjmrNKYCnQ71qeWF9W0LT/b9
j3Hi4OTm0uqmhAW3ffZMKjL7LSpHe3GqitPKhq/M4afYiajQAR/EvELL3kwkesWv/4H9hfKkUxpk
oHTQ38ko0MGAuNbIoojyviF9omO+dJuzKepEFPehJWBrEVZCIUAIzsu1K/5Ft7zZwD4CesUIGM7N
O/T3ZDMp2uxVbgwhV4PdQADK0j89lzin5dwHVx83vh2WvD1CD3ZQHn87tCSh318KnnSVCQHo8Y1x
u+pxHsTcN9FTv6/zHehtbaBd3sjam+Rj3hvfnI+tKy48J5nDLlm+hdxoNmZ4w04CNylzG4oNPZ+d
mIZexW3dDs8FpwF5yPn1z5F7dx8L5m9xXlRDs1/mmiiD05579cVscyn1LI8iwIi/gnXCCVWuapXA
VgZt5dxI8MSGfuLD6j9kvsHJMFaaEEKbfR5Ml5QFDJGYRb4aI7JS6OBA0lLX6WwGcwY7WbA6Y9SJ
YSPOexrR7r8B3zEXgdZvVF+nBUJuATWtGjy33fXN1ij2eCoFWxfENqHJ1pVVRFX0KeuWqy7GFtGP
v+9SkHUWO2IN76k2wOiyv7xoezBH7IMZN9/ZHoKrCVJtpifX+8LLZw28UJpNEmPVcn04gJZZDmsJ
CEPLsSGCQhfJjiHZ1mH0nRYy5bFcXI1SL+OG0pNGWxnSlEZjb2YS82pDNkq1wNeHJmDbsS72sT+6
lmwc7Upt9fpqlkkZYmRtMbdBa4f3B4RM+pXxHWaaieN4yqzsDJFJf7BxD6gGiEutK9reZNSbRY1L
3R1Z3GxXv+twqTncc7Bb39qPDNHZfHe2m7CNIcPMEjDBYvF+Kfbpk9oGbqADvIJTTcmjTiZXOQjp
pmIzQgNetMlZsYEPsGx8m/jgNvBvGNl3dtbEAS27WxEtMnMjqWn+YSZCOqUJxNe8H23lwtIhGCKp
6R9TbMzNBPenzqQSIYUVXOMypqUPDF9JmFj0Ehe6ZUjY66ftX30hb3OiX6z52x7kSJSGpl4qGo9f
PkfsYkLIhLPK56nvxih8ouZ1HptiJK54dka5GR6dC0prvrhyhO8ea1oKFo2qBUc4TkiMrGeMf2DF
kR4l22Pn7j1+/LBzQt+t2B/yfHk43dfDPFkEBqVotOUCawra5ZEc7deNlZ2S4vRLwPznNL9aTmTv
f8JFysfeFkYVtZfbyFYv6khnaOkzkTOiV2NyyQFGuj8eJfy+cu0+plLaE3nchSGLzbrPKCfjrptT
HWSiOVK4RhLhe6Ex3NzNcy0L0KhSkeg8477zm2Vt86/drnqfD6G2s7c1iVwgm5uSvazndjE3M4Sg
rFp7vJy4cjhGFKYQ/lA3rW74Z4Qf7ed91KheRei8nQYHqSgbsNU2enH8INOpMnM36JMHK6gYROlJ
TTFBffI36E85fb9gua6CTjP1tGkBlH415HqHCgZuDXATg/GUxECQRqAzi/yYvoHOWJ+sli9QtXcS
s5apTg73dIC+a3I/Ft5e091R8WKx3Hgr81oFXqJcK3HTEg5ylEIzPoM6i0PVf3vesap8u+gUU1Uq
N5tHXTW6qotY9+6cGSuM6YHruF6fpVxoEKUCf1CHffm0mglhLCOWQ05DK9pW6jo6TZmkQNotTBK4
72y0pBvCIkB37HD4x1xplAkz5WKkLRvFAv2Lpj7Wlz1gRbjJIp/fJZVsgol1qgUIaN8BSrjqYs4s
ynq5BD3oAr8D2EHlF0QyMdgmdxTr5BEZoIXyn5z75SkjrPgvqLjM9PbwzGk25FQFV85av6MwG2Su
7kQH3AwjHQ/Nstd+YZo09ka9PxAuPt5mp5zLOLQEuomH5/pylXuyxasI+vhEvVlix27PLybU+xpi
WDrrV8h/Uw9plDj9ylbLvcJx1JrchMVrurriBKf8iwYxnn+Ee3VX7DJDKsDNQ9ufIzto3kq51M17
wyKmSEQ3BRaU+eXWYRX/aFRRQskZhvL2V+5IfhueMkOIfvQstiT9YQ6KoebDDTghanbgokshZOBj
unsk17svW1GfpdgIyRRqWzuq6fsEdeJFjHtQMpcEhYSPwfzBBv5CnVIHfZiHbewJjikAyKSO4kgl
X069dsZZLiuB6W7/Wg1RDMAqcluN/7ib8JakQD2RvAf0rVzoWH6D4iQifwgOg+O5n+Fv5TqS7fUS
sZAPrwWInMJUBfnHGsk/m2rqsBWqx885xhzmapGmIdNAH5zD/WqAsrzDuWtNGIanxYQ3opYuuZ+g
rsFUnsHA4p3/Tl57V7vUDg/BHlW8cGiBGdJgIy0vt27I19SI/1Uh42pFLUrfvUUt1/jKJvRCppKg
QJg21dQl2HDz2tsribgZTaWZpBb9ZHtHz+oXvEMwyISk59tLfiX7vL4/c3AuAO/su2d4eufkKh1S
/JnVYQJM/snwx1c5lvXh5iFcnlBIvfYIbVyBw0rsRiaUYcZtVIi+rTqLmK4rhDQmZTfZBYKMGoKC
JCY0N4b4KcgP389Y/6ZnoamkDPhkuw03M3rjoFIvfnipwY2C/m+9js76RwgdM2G7T1RaZ02Kw+h+
dkZf/zaAn1fY+YI4ydD1CUqAiOEaTbuk04MK2IirZMqtyu2rPqcwD6VM7Wlf1l4imqdlT+bBGeTZ
21wi5U4OIUc96/SMEOUDEuvlXdsgNfH+u/R2rRHF8r21Z3b9x84veRhHC3mIC+MwXkDKa4jYKEa6
/eS6MNQ7Fb/m7z+glxLQakwtZcZoBpvTCMeU17rfTXfs3auVkEBw7Jb53QsJoq8vPcxvbQkZnAYG
lwveV6l55s+pDNlLduShhY7MQtnByvl5rckRxDcEv/QPlg60GZEGYp843oIoowBnG04Rd1pQaOwI
BtGg7tD7XHoOKS240SyOPTG3W4yFTzbrNq4kJnb8w3JhjKo4oe6bu4d+BJDkGEh4iQmNfzsjuWi7
ZadG3lvp95cvGZ/FJt1JQvj5026giDKCeJXgrCKi+ttaWPy2IgLL7tIaGo+C33bxRHS1t4q3LkFg
8AAdkQ51BVMiUhCM6ajY3Uw1kX6loQHJHsCU7DMVWX0VFi2TpQucrxkPO6sNyt6+uJnO/upedTZR
QK6KHgDGU0kBf3XBE2a918DoWRBIUttjn4B5lUgt3aqrQz5mpkJwMs5SWhlbj7C4HFQS4t4+ZjZC
YgGE8tVgcjUVKKEw9DpRXVlXvt4hFPXQMt+YJZEW3vDwzV6OPukU/s5gvXekREgWL4mfD0SF15N1
BomPMZo7j3IDXhYEIu91j0lbVTCc1c1T9nDi+CJ3BZRxLg5BVm3xoXjpJFgLRUzHamEZOzeC+OEY
mLEzjRAvo+/PJ2+gCBMYK3w27Rtf/yMwfl2tbvt8JwE9o5wcX5IXk89AmF36BFzj5XUFy4r+2yER
bT3DyShc7r3NzEbOiHVvSLPEiStSEpMSvDUY59JHccEi00ejSKIaw2gZrRwq52J13/GZ4a31QxOy
TDrV6C+n8kpsI3F6Bp/02qCWUFTgoxj8WRGZjrhWThZznfOdr9YvvFAUpAUh9Q55KdvYb1vKGIJ3
2XzYZt1yJ19lUxHsoJ0iRhF33kCKrnHQgZ0KuBi3kKFJO4ix8iLCKvIRFqZT0DjZt/WlB/9cSbry
4XEDBHlvy2sL6mGu1TEdwo+Xj5Rw94twktg0fLnFH4E1HXwi1gZNZCqBGjqtS2dkVCzHdf+2LqTf
0d+hxZ8SGjOZ507FS75ocGVHKPJFUfL2Xw1znbtqBV6x9P0tbHLKeNVrn39Cg1NWGaDM7Deh8RSh
GZWrhjg0bIEbsHMBENCguhi5x4sa/MM2kSrjSVv3RNgki5jvrb9A/tEulNwtuEObgHS6iI9r1JC0
P8SN/Tfr5ZBazk0exgILYwGH+AauDYe90Dm4ZlaYHDx3pWFxEaAbjedtmzKuhdK8Ah8ZSS6NghYx
WQmLe8rZQR/kRGhBOEjhGR+Vhg9G51fMoElwWfVWAuCtfz9kAkfjPYWTKaojoxCqZqbHce8XSa82
49Bq3w66Sflpo1Kh68Ss9e4+VGwng7SRBZLXdQef6xVmVZNpjSriGf8VcKWmtCagFvXXdG61FiAM
3KeZItzveCkhJ2UEC7zgtu6cJpnJaQauNBG05Sl8qRQSYNn6KY+ECuKHfgpFlrYRZqiYDEV/BvQP
yIcNWACmU9dmpWmQ3tRX1YrulfNRmNuVxTLwDTwhHW9PyFHlTK3tXAcV7X9SadLnMkIhz35GUT+Z
hU8aJLxA5WfhAYVrAM6QPnhvwOxk3Ry5goteJvthFZEVVB5HKy16NB/6PODSNftsH2FCFb2uieFZ
qknoJWES/w7GzijSux1S03lx7wdMON5U+2Yqrttpq0uYOjqYXb6nb3Mayxa5IWwoDQ+NFM0snExk
uX/6Te9j0tW8GWZYnrKY62j3heCKN6Qsv2ULkJoqKr9X5ScOBtofVmxeJu1W3MxFoKEKDjSgTYZX
3MS0qK/SA9l3GPwClqtXvXHTQxNnFsj29FFQmvA2R2OTK+JgWH+MZZgjVPZenb0mThvecXaYUs9V
rWhDfdEv1VBnjZ1k/tNUHUNms1VM9h50aV34hX0zOu+Y47xRqdG+FIhUqqp0Twzas0zrmneRi6i5
zy5GBLZTe3ixxwTLomDxFjYHR486IDrB2mZvREqVr26P/P4QFY7qf3stsbeVo9J+sDUqaDCO67oS
0QlRSfyDWk5wCDZsiT8IljuY0fKEaqNLaPC/pYxrplw9JntDNVmfe+aa4Y9/joEUI0nOLU6Wvz+g
efPo8HM04oJwuZ1NDi2eU5VEMTc6wllvOm3kqDo/agyhzTUvsJF95IFqLsXGH/p8wcyEMiy4eOo4
a2sAArwQUWaWLbzG6SS1WC7LNWUCEMwGRzmTduKk3/eFKKxQmYzRAs2019YR1UGsHJstFx9hro8I
8iADGTmXUEtuSGXoOHp9vnZlO9qkK1fHBNzIOtNlAjlXk47lW9sAvT5lw3vZA84vGNv9oQh0fgcL
JZD5cNfswTQ5I0Me8S+QICPg+Lb3FND2pEwCde6l7cycL/vU7C7WSPL1InvjOn61cjewrwObzETX
sx24OqFuo3juscu0BqB/eAzbaxZuY2gOjtmOefLzzpdLoOkuHvweoNqPYSTziny/s9Qllm7ti7pK
DD1rHF8I8jcXRzvhyIZ8AghK+ZSal2xFyUYGU+ua77IAe0jsW0FPtSecj4UZfz8qEQbXP7CCBh0i
dlb4y2/sCa4+mTqsHFHowlyM+qaaGJtawsRAYwizxpfY9pBIQde1uNxji3cojCcCQphKrwOnbL12
8B0PtglGLohr/R/3SiGTanxlZpGEGspl/IcpSLogD9zkveu5M0QUWmv0cXXpXHrfvGd0x/XYRNlN
wHKVPxOc5Qg1/gjlL0JHMzYUlqW+57rXC0A6+QtmYnlRN5UxCGycfJFRf/NDNbSKS0STHUEYgh9t
s03vsfNO+0+HPEHBHf45K0v1kyn82saK2Hcqsy5/jwtMkPeyN3Q5ekUGB0VFHLXXOi9gr2xlNcmi
4jxde3J/xbtS/km8ncq5kQMVFlIc+jTyRn3aHv8Md+7qfaSTb/DvR+HL7s3Xk24g3MO4dnE/nfrq
El9QbBFQnBT67lp7bwgZ9/wxnT2OCRI8IDWINVqzInOyRbYDFfS6pJg9//MSIDx84ptKTwmglKqD
/13Ow+NOgdjmZDhdV1jc0EQ03JNv/K3Eytt1f/ujjQnAKpH7Pt7a6EUEyChU5a9Vcp256gW7tvxp
q20J9duOmvLm31DNczuish75h2v3Rq+2QB/G7pMxcXUvxeDJT+L//5kneJSfzDYGEeXnJbn7u2zE
5NUii/EaACaf0j3tu1kidSezRt8mkzwFf6UgMmWNkSZQ4CWcvGdQRzMzJKLb0qQNDfWmz+mOgnyI
cUQBaFNd9K2xuMH5mp66ZmJrWcimIn9TPbCfwBBfGl3TDwqOrOtRCS8ihAklXNk/jYRVql1rPIjW
FPeQ7mHo4DCzhWNfXLOnEL83FMhPOtLJCKkoOtL/zq+tI0zlMd3fEKGb+qPV1hvfblFgQ13OaP0Y
BaawuY+0NwGnrACRPRtS885hnvFM58pvSGR5GgBMj7871QQfw/Kn89NBRSPveqB0D8QA3pZu1Z/i
MzIj8E9B+u2m0ALm1ftAvHgyuCjGzANdtt8SYfv6Rk4iyJNFHrAso0jpkoC21WmYhC3MNsyCpZZZ
AbzyqkJVYA4tja0sxnc+cwxzYF+Jd74z/oxwHOZghGa4jXuq8Qrt0mjiFx1hDD9G88QPgL1RJm+0
zEi8MfS9PEiFRaq4YwwuEW4Du68wlwOd7TRujSX9FXm48ok8zqMuxbuXzv4S4J+Wsm8KZOKkBCiw
KLnzVz26o1r10NQJfeErNuQRLTY25p8WnLHC6lCO5Z9F2Bul6U7RB8yj3j2nNaUWR1KAY3CSwHPA
ndGtTnyVxy3J0Q0mh3oq0499E/pzG8cFCY9GJKM/svfnRP4E9o6irVgmWKyokEp76mzTCdY6MvcC
tzN1o0UrRCuCIMMcca29jaS1d7k1FpRzS/Wn1NAwix62G37dcRVb+25O6fKcqHg44SixwVji+F4K
PQo5yuWC5ewxXYql5wNqfL/So7AbbJ3tAQXthRAYcknGUuT5+v4XM5uDFtztKd4w6Xv5Ymj0rTr6
FelPOc/zmLT1eaSaw+6GF8Lw6+lLnX3BeKvCOjKJovD2SbyQXImv1EQ0oVEsam++4ZYAoW5oie67
fZVw2i/G9mVTdT5Y0TssRpS++g3SNAGNtBUSuEBJhdNE6yCXEEHMIcoLD8RB5ST36r/F921itDHz
cWZUDHn/nEu+S+n8kZr5TbqREjmhsMINKsM2MTB4RkWGSsOuUzDFalzXsnaBOkctjiKMTbP8SK9I
/eJs7J+8WnBKQ9e4gImU+F03b2RAXHLQ/bJDVKXzZe0I21qYWvr52GIuqO1KkAD4YHP/sN67qKbP
zBTAd7Hf/jayVUP8yiVy8pRN9gPTS5H4ixNU7ODJkPJ9FH6jQpK2AO+cQts1IQPwrSIbuRgzeEJc
ECaZev8GenPtv7p2Eg0xExc8vg/dZGGKVB1vnf95dr9BTVJwifHrDQVnSYGNV0AK5sZqPW6gb7mY
2ZxFh1tAt3TF/IUkCTK0Qr69TmPIiKGqhOMBp6tLK31b2Z22cyJvNzQEdtRKhf3L0E9FU6ljA9vm
WaKf3ULS3lZgvLveMrv05l3TP2e/hPjCz8R7+0GARKwr5AFtaAsRJ32H8NGxgNd49JFK9G7wYb3U
RZCfG1FdBEXxWobq+y6K4HFpwWy0Ll/VUEwvWBngxaNJwapXWD2mi5nR5wKb6GE+qsZxdfmPvKbI
AJNPX7Lw9QTzUe98+A7jwEpraGR5hwV7i33jrpUvq0un0K8w3HNUh19mH4O+Oi59irJ2T8yDUj+0
/mgmHmlWW+NXBCV+Fse/CkWSfZmlnQvRmecYpHwN/vC9IzU5WR682HB372yMUyxMekakqZYXuM/C
65nWa8c0VxGAscF96sdMraHR+1Oic6UMXFvZWA8b6DlWKpdirWSP00Kt+iAfrpWHIablelrPLM5I
xq9IlYhSCSfMqpG9SIVfC0fpkY+D2+812jTitkIIEodOVBsJC6j+3mJSXouDpe1h4mPktpzcL8sH
ocDPZYhoECzRGKZVSQT8KIlcLNUWpQsOUKnvEnKWH6w4fKpVP32mVFzV2bi4fOqbQFAtYa6gzfra
DOUMb9CQEYr2pYnXX3j/jDlC6ucv68pPt/QFYj2iNSs8ffrGZND1WwS/n1ZSPA9uykww+oZ3PzSR
fKNAzLPk+15jC01f2rFcG8DEclYvSMR0wsvRQXOwuPKSkB/06XGkBSUDxseh+xLJq1UYbq3vNDdq
9mKPUvRuFZMzKdqe827e7J3fk7ltD/a3nHBdGE1qFeuBHc9F2T8iYUjCRUq39yMIz1KQzJQgdJKq
nFzEwNeHD0UYoDQ3Cc5g7cJae3bNSZG/nHUP5UkUoCUTB1OppWT51BV+tCyUfA1vwiAXy5I+W+ZY
kWhXdUWA7rgcvsSTRV680rNENPBlWtt9zcrF3MzeHQSZGk3mG8P96GytGG9ZhGJPSZjFHVeVBad9
NOn+5ETA4ZGf24+OyAMRHmr3RibCw8c71stS8RqanyaH7EEY8LzrEca5nObSdj3LSv2VEXNuPaX8
qp0QOfKGpUkaZWp91d94oRSrNLpDQwI7B0rwm+C46QmUINC78xwPvVoacmKCR0Taa/S0saBkBOfI
Ijqn71xxcu6EDpbbkCj/UV+jka21SeQv9Mn5/TFNK5NDKky86pA83xdm95WiFQ8NG4iXcvuMlbuU
RdTrtqrpZunrYBvX4fInIE/Q635PC0S+lIidDdYsCQ/iiOQL986JT2Y/CDccWZriytvEgb/+21vo
1pTGLOWCaNBQUc5iBxt025G5q5ajGK1P5oyqb049CQgoqqbeOgDSpil6XRoacQJp8SeLiLUkuJnb
PpUUIRSqE1k2d4oGiSMrQsQVTuTwi+Xyq0HG3okKGM1osEaKGjpUzJigKygNTiVqv1Zyu/RhRCPZ
QqvNUY/fTqR5oHi2fF/a4BTyiiKXOUY6NP3ZhYTGPhjEqdbEkIXQY9jsm3LE7TmbN3O0zEIBP/uy
GyWWyNni3HtiCIQzguZ1UOBxdpADWZEuk1q5bua4cFbnfbsknLXZCJTYWFK+Crh/tklH6yli3Fhe
LHf4F86f+tzk2Yps6FYQpY5aRFbFP0tECpVIxzYK6cfX7zjdmAPzZ0tXzwY9O04gcowZzIS3d0Dw
Wg6siXPuzjZDL7M3RrHZoSiF3wU14kYW6bnLdDz3aqU+d8SEe0mQmykjrugmEl8Ji/YAi9uuYcDa
lGbKSHuLKyr90Zzc5/CeurB4AY+mz6/0LZlGQWBAMUf3udSGMKMYNBCoSaorEnPVqgZSeGQ23KyE
cvHdILleMu1FEwZ5ayeUVPScyA5+aD2RMMRRd5jo2ku7ey0tptZ2Um5qWhsF9S3eKRpiOhz/HKYL
dPTfoP08p1ZsN6mXFOuhS+zgUXOKJbyuyq3qU/MIKbSoak+aZ/7dB1OZbyCGX0Z1igtA9NL3K+dw
wPdseJeeRGQrPmbsS83oWu0L0ZrACRgo0lNVbxzHugwbFdjeteBcjc1pZREZLQXCw3mZKKGyliQg
WGhQj17N4uVsNaoYQ44Z0qkFcct244ytoIJ0Cc3nQhm11V0s7j45lyA0hPWsQJP8XwlW68Bn/42J
j4ABzrZnQVvH2Qc0Hdf6VU4xVyhp4flfE92omht7cRJfVTrfSMVk7blES8JLXZH51aj+VwrRQV/v
0GnLMubHWmFD6BrcQh00oPszJBppcStWSMu3okuPyFTqqyvFS1kS2uFDC1KBqRtt8plaAXnlD2yZ
IBiU6TPtwSUEpgSlnbnRmnFOKdpStIj/5k+H9tdwZXfvZrF6sk2DfgDYSkdvqGr1JTrsKMRsd1Ti
PVTteSRPulWEP+CYK1H+pCz4hTBwwCSTE/ciheXcTEywhVR9nyRXoQZcfPtSIM9ENvfdmrcNCu2A
tQ++G1UgideCd+NvkxX4zdsFLlyR050k//15TsbEcC7T59241nCKpaXr7as766ojb8F5BujQ/ZXK
7ZyfXSPiqvkn8C27mxDxbIHU0v9HPSe5sZPnhJbjJCWkC4eMsnvNTO27JILxxpWOpsWdUMTygKSR
Ato3Qm4gFvHF5ZFeoG5S82qcEs1f49d1rgI6DdFCLjg677DiEN1CEn582y0OEJeRvZspMgjLoSsa
ngiFnoBZnnFtrkf8qSfHMlB3IM+Cu0ku5cXnBJdDci9llPXsb/cVpH7B9uV3uzyiEFE6Vy2ypvv7
yFFMA7A+pVrcy6+eb2JDwKXd9TiU3YBR2YGy62RH5NnSl2QNUa6gDJ+EYzfIlgTM3zu0ptepFHsu
o/sMR/NmbVa5EbVuEHOFHpU4UkwQ7e7efv5KIgb2CWeA80YDLdGXifo8WaAarXbpZOP5nCuN1syy
cYHNUHaE0vh10KKyCEfzHSssefjJEkqbRetrf/fLQ7hA09vou6GAgM31l3qlnn5K3XVwtzk8TxYa
Z3Vdl9u91ehR4i2sjjfQvPC1p5lvVnjyK2OEHMeVRk9S18uQvoxWXdI2vtpv/n4HiVopSBf2iCQQ
EGTXMdIEnf7GAa0/Qf5bHVgemPa7hdN0LCEwcz4iP5UwEV88D02OVVSd+h0494rHILx7O8YjHVDi
SvgA4dn02HMVsd41Yx55PXbzMFuqNsDK4eLbMm3MxeHMmCAMOOOwzJ81WFXuGKEhnKHFyl/WUOnT
I3PFAgNL8Ri/e2R0sHXaXNNrxisu/LbvVd2yyGWRmR+avLKEF4cAfSuMYTw++PYTbPZFfQzc0Weg
9sw0+n2z+9osXcL7joBqdd4xP1x9ow2UbQG9Mj/vUYxGhCsiyXTQOI14DlovKnLEH2fPhbblZKWq
F7TBhSy9AffGZjqn42NvcEp4+mBQaxuIuLH6Yuxa9Rj0nm40+8EDxTmLpebGLVbLgGya8QblclBe
0DxoaziYEMkIxnNKPVpDzBIOvOuIHdgyt86KPhRcO7iglQe7G9x5lvPeU2i3uuc3TQgt/U6U1Dt/
X3PND640O+Iw3i+DvCV7yvDqBU72YwujAfRChkKMPJArsNVgpri9Fhwlz/21mWiWgeZH7XaEmy3R
d614J5cJQ1fC3S9QAtczJljuJYlc1uLgOEPfSCDF7pJjTRQvlrr486AMFNhgYr2qTta/FM+qnLJv
/uv9EwtrMWDtQgp67XV/p/TuE5JHilfXCQSoLwWNbALw3N69EmTbcx791We+DaWKkndocYSuHoVL
9Bu8XI1A6G7GBxiFIz2VfcxDtSL+V7GUbqh6SA7fHQB++zGpX3lAbXVFS5KXn1J+qs9ELd3N9QJe
4eJJxdj8whFVFaLEg5stMsHz7U/R1V3vZh3bI9hLM/d9jaGBOKC6wXRk0mVr+VzuvvwhKeJryJt7
PSvKSx3abFoz97oBpLIkhvcAn41bx+gPPjIlxxDY6l3eey+CWpScGezopZaWcHuiqSK7G2C+lFG2
lW0U7n/ItuN2OVBLGhaeUFMahuPeaXpveRRe9T/c6LuQEEmJT6TmWVqSzR4kCwszOKIy+FsDOn49
stcdQjsdsXcKnZFw3/uAQR5mmqgDCgupUwiCK5QQdTy9js69AU673zKOtIria75TvAe5acI6SmLk
n941ZgVVbHAMuB2JI3TNQQ761JFyBhvhQ74oDGL3wxd/OpLfJ9/apuKSjej+TBGxpZ2HV/f+sU3Y
L65MkGGLqeb7DoQ8ieh90L+VnuE0RlUV6rt7fX7tCXz7vO66BcmjHjb0p4cEigE7wyz3TaY+HJb4
Ktvh923GSbvCmH1VNSJIEIPD91rvNlgeo8SSyiS78viqdcD8SlrrckiwEBlXflBPZzu9yCct1f6R
cka4JtetDj1No8o6HT9TUp1eiDA4vv/iJAUp9jo7SM8VsmaEehdFgyj8vbpCvGhb14ymp2Hm/eq+
VG8JJ/yC6QdiWddaYtEBfUIlungoauw5WiV1Lt2asFGBxP2XXezG6ZSB/Uzdzj1oeL20+I6AQflZ
UDZZRrKsZMlGac42eAQjDaHLIushSTTC6WIDLO4w5Ewwzo01BXry7fx0bEgcZApO0tuQ1Hw5sXDP
oiMGo6fAV+SH02Tr9q2tllJW+AbtXADjNDl5s3GgCIzxt1+h13kqbOi6BSXeRluMqLHT7EUes2zn
nSB88hIQfm45otZdhY5Oqj5oLkwaPXqEa7JNtx5N/dhcWhKqtxfDAV2RypHtXYFDmZXf8spxe8fd
xl3ma+rRpo3VRRch9CHzGxRaTZ1t7t9+8n0qMzAT9YLJkjl3vWcteq0vHw6qN/+x2guBcKSovF8F
7FEuVnyZHAtfsdp0Lomks2+N1nt7txCqZ2dyI/bJCFIOcPSAeuu5M9X6brrAJA1Yi/0upMv76cz4
EVGkoVVS0HmsLxKF/ND9LUXK359uUhTVtuColbBESU3SaON8HuxmaSx17i+twA3eaGsGmTVJ9H2I
Pnz5kTqmsVKNgY//K2ZAb40dmnP9Ma3gLb9PdC/zDklyBF+IB829kffqgPslw8auvxzjQqTva7C+
IK5bsN4UQn3c5/GipRrQ5Q96hvYDQPYNa+SX6WDqqGOP1j/J3Cx1kjtZuEZea3U64RhudKcogaM3
1vVPXlR8U1VgIy90/iZMujQQPCH+cRBOOXQhgNGLpfK3/0xDAJxF5Sdi/56AFy2zlxCYh/8iqHZY
iphPH8Ut7EzKnU0jzhK9pOKt+DlTTnTtWGbggJkq8xAjdu79YbQ/5NwqsV/laKak3E/DU42PBGbe
mEtI89KKle1zyGa9nhobI4PoOeHxFJcTeYe2F4sJwrXQRwVobcjmIYhJTkoxKXnarVMuFSJF9GR0
7MMpNG65e8zTwGBNIIzxASn8sIW7RoyWGE0n4lIVr8wmbuxgrvl50vm/OF7e+9O3jq0UBV6G7gBi
mDOsVRaT5OybaTHDb5AHHUIYrOK8LnOpx7TR+k8mrQyhBLj3mSLA2I+lA3LoFBRst+tCdZNE642f
8GYuIUl4T46q5HSXlkhqYDDrpNloGPOR8Mf0d/ygvX5TZP+4HwwKZCg7YKOIvyCzHRrpP1mmN1SU
4KSbiRJPuybToLLnkvi27Q7pLnAezRGlQdfaFNU5pGZpFZrY3PBP9sjbqdhUe+BQlCQB/xMob1sW
JV+sqKwvhl6QoaRFQHo7aKyDbPoOvNG6jdjXYph7CNyxzunXrRGqd5FQDxGuZpLW7Vhogh+chz42
rk1HysNK564Pn6m6/vFF8v7Fm790ukcHfc5gdT1SVlUyTVDq+M7MRgjzkxun+4LW5Ag6bo60ApUr
LtJC1ywKdToQpOkSIXGY/NuJ/Rsy5CdhRAhbd8lbu+ttOjRgf+yyA229f3gFtfPQzSkE8dgrXPaf
+eocBV9lLnbbZ4A+11u6Q3TNCdVxnSqX1HK2RNwfbLbZ/oTq4EyNRDWoivdXq2OuDtmOglTFAyXS
MYCrqfy1X7v/JeZb9qQQHBd7no57l9zwkJZHVnmKve3dyNnI+sWRx7izoQMdXujCG4odWPjX1Kqv
gewhopMHBwH5/5DJWmyKDyoVIt41wL4x53Kxo27wjnYRafEXYSQqn1+ziFTpigFr343G3OxQMrpS
09DltThviilhoAWIi+j9D5LRt5mNv+qBTR+n8190s/MPvV4v0NGoQZWdy+8dcZG0zSz+KzqpCphM
HJKpwtBOeQTRisAoT9gTJw3HRu9tixbdrvzuEUzEepq916exVR9B7l++vlfa3GDNQ8CvdgY8SWp6
CiHn753POHBdV5Y7mM9nEYABQBmNqSReCRKeZp17k9hecKcTcae0UraaPxArLtFPGxPmB9lW6Q9u
dS74lp9Et8kMzdQHtpVE/fW94afA5WdzoVFScq2AHvqarfbknyb365unx7CHAQ57H+CIPJucsz0G
rRdBr80VQL3EX5xYIjUwJNxgyPdVcoBsNj5nJ4npV5h2HoPadHNFyvzAJYXnLIRJlzA4XdSiKr40
CegaVIjye5UdSWXcw22sNyUHgLJaTUzpv6W6u/lYWgxuaSpB8nyetz3Z8qxevoB84F+hoH6AwIrv
eVgQAlFeUUU8vK7F/SDGb0VA1zJw2aYGVs9IzhQDHDJjQNvkJFZ2grk8XTUwINBg5njsomHgs9Po
Fu11+4V1O8DEdC5DPEBEXs4DGH0MiAT6Aazj7b3flEFC9GP6LnetqFgtrDqohfBhJC0eX4i94BUm
NLL0kYDrVP6wkKwX8DB8GGlb9n68SUIrKBQjbxqXPJB7CP139DpRYosnJYOzAD5DKCTH6t9f1Qus
pP5R3G6fPapVytP3qCFhXCL6sxXc/QncNWcLf4gIhARsCUQxc03k1evLaMjsaEiu1+TcHUmdqW0M
g+fUo4I+e4mEvvy425Zl8NhgIpst5+dNJzro6eZaCfKzKjGCnS6w6K6M5nPi7WgzzFSDXaP/e3fd
W2qcQvirhYFxxOWxicWXzvnUyIpfXMkEIW5kt6vg+wZ/NdyVPq9pTgouEGbz7vBPN/B0h3fL+mT3
WPelIfr5yzg0VqNXK7K3MoNw/rRQD6JPE3EbMAvj2/i5MMLp5gJQbnXdKPFbBoSAKz1OjvbLZ62v
aVz8ZwFG0sUxOKv0mtNPKUiZpQ8JQn3/NdFcgB5Lz05HgDl+BPNtXWs4Yk2QIWtJNM+hc0gtP0pk
p3L/x4yUe+POxFIQMd42QEXWqMg5JE8YDgud0pi4Tn0z+dN6hVB3eS6cl46Sucm9/Xm5InFyZHa5
9VwmhaILmLGR+AqHKzqPV0HXsb4O6TiTAdVRQpharLi/ZMVVQBucwXD/gCuUA6b9IXqKmiAtFiKt
9fBLDzQd3nQZ99xdlt2QXNKHuccVBc4S104JLwPfcCerIAVXsxwk6JWv8E/ncJaIAfl3iNQD3Xf0
6yb0WwbXIO4urun5xrgJpNsZ/iqWo3J2AbIi2f30/Sj0Q55/nNG6vp1tGsHb/hQqB2B0uBCczV8u
kG6HPGZ7JJllQaVRo2r1jV6Mc4cKTG7HA9eUFdSAJbptG/HKBOK0uIvzZlAPTaOt4siDsMm4N4ES
lmGv8i7GBPEjjNjE7SIrXRopEpkasGWoHXUijryBfmDlg/1QGtjK3/RjG2Q4m34tnvSEv6mcwZnR
YcQM93ooRkFTctyp4TBRkXqmVu40efmEwPH7A+N4cUkg4Ki2V/26s3V0y9QEyzQDhKB5JLJ91jor
0rtmbAHqcxqhaRGUGT+e05cbr7O0fA5vyWiccwS9n/VZJ3PnKgFRG9j8cl75WXmeUoMFxaiAENJT
l7nNRK0ozeDZ9PCp1W9HjNibaswM2Iyxj3hZHDTnJblkgEga8/OZsjj1JCmfKosflkcPdowCIFf3
FbdS3YXh4hqz+q7qjKuN8cLXTgT9xWtdT83PrAPtgGir8/dwEYw4QBIf7EwvimNRSJunKaIcbh6J
cV1PjnXQ2iudSiNWyB7eUuwc/Jt5zrmoDNKH/nJgBVKsBTP6MdsGRbLTHSu5EWhZCKeW443D8g8A
CxXi4jrIjbHmxJESRvwIz9McZMgxNGI7G1/QW0VEs8/WAEgqNBfer2ZqSz93kLoIJV9sqf/r5bke
2k0YrdhiZmARI148kHXmzRdOtqVMnahWvWGiSlOTu2yqCQEcedFmF/V0Sc2bRmCuxQ8Z5n3VLW2Z
+xSQta+amuFFLb/htZpvbqL+eYqUoNP+fkmLe8vQ5n6z8OaS535z1mXHqseO0tw7NpV+/Wlb06cN
GGY3R/7pFU/8XD/nshtORBzdDXhNDAJ0kdhzYkbyVGE27QKAO2H0ccTqvtAMemRcz+SyDDUkjAB9
RD8+jnWBfJnVjxoOL6Tqg0YFonNKgzwuW45fRSzBe8TP8WG/1NzmIx+ux9oXvkySSPPnCd21dUdY
MzxdrJPiJ75ZsjSIrh9aTAp19R4ArwRlCMUipcF1RnPoiAkCKIjJdRuR2t7Kxa3ABKE0T82vzfCX
NhxJ61cABd97koBdDg80pnZKEU4FNmviHSHDghoEv04y5dDh03ck3vTXc4RXLX5gaFuSm3MzkNdf
EqePRWcXrOVw+BRXSoiezpwQi0Pg7TXc8mqNsnsGDJ3/tJGltx5IS5lbiyaDLjzlNNSBZliFpmvL
zBpLAQbmS4KU/0qH6GbIORjEZZTza3rcc6ZqkpkJ/dhVC1mXGIVosQXnWkAdwwZiv4rSJgtACZMQ
19ob3yj15htIygsZj8vqa1an7nxsz3lqU+gkF4IdtuXWTQrMb45VzSNB9UOWCRrogADpdWw3C71M
NaXZFVDDmmc90J/gPDZD3DLJ/N/5mzS4w9nhRGQMtNivu7/eCD4Fecld7Nx5wD8j/R+h5jICK8F5
2KA+vbEkZ98GRfJfUm0Bt4JYARhIHy1N5E1ElGDeO+091PeELq/bX5Jog9pfWmM+ZjuK+d+dy4Pd
Dt6Fg3SXxip5xAyUkiOQddpMIqS+SxGJhJswcJKvHYLZ8DKmNFj07Hu1jzKDLX/Id+IIcRO4bGJI
tfVz38VBGtqNeF7UcFkp8N/aJd+Q0vqkAlcLt7uNhB5tNrPobycwuFCRL/YTFQRUgduPosaMYMuY
QL+FRihgrQrZmsy4yYXbs+QOz9Oz44cnPNLyUmfGFzyd4YMgqVIkVBmHvjaiYj56E9mwpmCI76bN
iJrQEvXPzgoXMthswWrHD+gzexLnFb+KvggJfz1hIk0xAi1mqwoXQlK8SSMXbgbfw+BloRYwymC7
a3jSx1tl7ik1Jp3AlSPVrGLWPYMp/rjbYIz9msAZh005lRtB4zRfm/ppVX22UuWuCtC2MVCuug19
YhqF2F8eBDiMYESzJoOUSllqnL9oZY2rpbKyXLDQ0Ij/Akc85x3s36nrDRhD0GMm8PJlkBUGnHLL
1h//c4WERwQ0BmR69Hz3vRhfXPM3Vld7rP7nEw4chGoistlWgFp7WTP5EGTngSnoFbuP6kD7QAFu
NZG9EHrF6TdN3ZNQUYU25hkRuBQWjlK/micaW1pSB0QpCzIe+tu+FVNn8nx2facSO14oUO2yaD9G
6BDjumSZrLYacW42r1bc2WJwLUjRsMB7nRSNEBWnqXoV1wQcvZBhnsE/aBThmRrSSgu8IO+xn4VG
w2JpOthqqbo57/xDgTQsleBaEBwbVoz6qaUzkaU4hP1lh7xx2VzxcBsR9MZYSF3beko4qZOMNaU5
7TZCCQ7kvw5WgKB8RbvdBhy4T6prU9OkWkxbvJviWBdQQ8oFZqv4Wc+gyIver6dZZ9oph15xGrbB
BaE99pLKB1kkFbXHk4FI1K5+l2ykwahpok9Cp+YPZ2UtFkRSRRHvJCIclNtyXg7wGEut+z4ii2yW
gyktG1U0w17UQXalydBiOhRaLQQStw20fAN1rUGw7WgCJ85xjKAPXPLmIgA4HoOHMx8DEssAJA8z
ClE8gxuD4OT/8u47C+w4nUn73dY478c+3sFcgDbVOhHmOJfs+J18Tp5OYRCK7mzcMPNVqnqn0MDE
GF2L4Og5j1C2c+6QiO1wxeBinR8Q++hIvs/r3jV8M9jfP6wVFYBYeCIsWv/mEwH2pffmAmLPkWce
GykMdRFSjLjzY7Pt7Ff5rnGZgJxe5CRDrKNhAwNBezTC8U29ruJh6vuGsxEt7LlGipQfNTE2VVky
QUBMq7EZHztNfGwQfrmSUxlMUNMB3OD/j72CBSnVRWjGh8VuL1Fu2x8DF6tzVNzOUAOn9eTuv6BN
bWo1u+Oj1PgiXckM8JEh/1EjW70B9rrfRVOdWcULY5H243vsJg6H/6snjFnO21CP3R/rD+PM6jgC
17P6YiOtQjyrmNw2SG2B7vyvKmK0rbFPJ+sCCf0DTmm2rVDsawbo3uBmrLNCG8DM+Krxq8Tr+qJa
GUIB02y7nk7m+DoBuGEFgEWTHsT75uRc/3hRzBrDVvwM+NNCI3w5TVfCjOnbPrki7dmEjU3MuBYu
Qj2xXRHyxZAHqkWIEoD6CyrDr1bx2AcaGZikT+tSnxSRdAjR61wi+SeJbP+7ckkKk5F+zCqz2zb+
B8VJcQP3OsaNmaJISioHNS72VIi9ji2yH2JNCiJGi6LoIZpS0vVvAvbK7rc68TkYxh1TyusrdMqZ
qm2khq1Ks8ClMR+b9VfCbGK4p5yXfbnTwPVWUp1UVtAfBn+cM4OUiLGZNKWFBeuaaLz2XThIyrKx
HVk1Dmvv37uFL6a7Oi0+KCEhiFgfBMwXapnnYL0dpKTRx9JayjJKlUkEWZOMocU2hwEwIAbFgqR2
oW0A2GiUdn8IZxUEJWo/MPm+fR6OP/cEffzaXEMtW0mXokLbVY8MSbWQgwPUpRxCjyPvwffTwOFC
N3X1YCIu+SnekMHHvoJTvXCKPObuspC5zguOhxlNwc2N9K4KiQPp2RmlPdeI5Da0jNs3zQtdxCX2
La4HEkQuJS6GtfQMN8bVHZvcJ2oOa0qUWpXub67XIgxMsEIejG0kECld29a2FKnVnToc9lYFlUhb
xWZFdimZSCgaXYUyBL/bHdlFWldgGmc/PeMKA6Lmm5s+oaGOVkFOGK94872i2vsF2VyeNMdcOdOJ
zBBb5QDWMjvE+p4qGbCGNyEKxHQke2fUaPGAiHgOiXCZXEpdv3Gd8+jTDmtRAKj+JG16VANjloDS
D5RfG2nGfSQZms3K0TE+qZQ61q/znzuTNoeNv4SuHJp79ou0eBXr2e4V+Fm6s+zbNsRhWyHo+AQG
yazaTfkEyoe0QYaZFL8Fgj7H5iYo1MidzELQECSqTQR2zULJ87s/0jWSt37njeYH4mAV23BaxKOG
M5O3qXjLtDGXP2lFkqow4Ccu9dsaEwZhtNRu49jjGp0R5+6t9aAOnyN1K+jdrpIjdEZq6AKko5nJ
rcXGDsT/MLT/XQTKWXbldUGXwyl+PLqCTqCosiUnZx1rKPQ1uNKgg1bFxM7hiwUnbPP8n7pZdCpm
uvKrMlm/2Sx06lWCLPVaD8Q6HRtqdythQ09MhfKfw1lWVCKVATK54XBEn/T8pmvLUA6Q9YNE+pvC
9pYXLGiGtsS2SH9efKRjhNF7VXo/ZksL8+xr/k/V9khZeDcEs6147oCPRU+O+QaIzlCXBFZ08zLL
TCC8loH0hxBAZN+xeuF1vNOMfQZ/YI8kNYN0oOo9+gbHM8y8bOVaEukm9ATjhMFyiyZ67HB4M0DL
KMj3YHUE1PyT4klh9TLPa5jZyEZTHVhxYIdG3CVVFrMQZScDFeJmp64q2a+GLoU2wlTdkJ/Q+S6c
ZlUhtH2bjqyD8uCnNSZrHGwYYzcQhxmTpdkdJtfle9hGEEzJMeAXLzy5KGl5ptavvDFB3CTILG93
K91GPhM58UJz2wjlD6Vkf1SQXPX74qA7BISvzFRHet5EPDRyWY80IDSejPrOzUEVM353opGm8FzB
kqUsoK2E7rXm8CP0s1F0lQVP+lhYro+bKbtOMU2PdRskCEbxlSOybrOhKrX6rA8/r8wS4hyjFDId
bCP66NDziyUIXiA2kn7G9AakMoeu5v9MWpigHUys60UA6ImGkmSPqYn9Fm9ODu2oaE+CT7nDQPxY
FLqVUjg9nMj2sER+FWMYlElR3hd9OBgSZ8ie4ApfDQa7b5ZNVn57F4R+xY3ESD/6tPQF0XsxEVGe
Oo6DbjMh3mwLJqODwAkQY10eOZL9GbbwQmhx1zpB7t8sfZWlBufMdsetwVf7vxX6Iockq3/pN49v
I6Y7E/SW2MwVF8b6WPhh0jZmUaoAYL+SYu4OSB0IaDP4z+kmzAYCIHVU7QN+H4ZGUXkas/hokmzj
keuSsA67qgFHSBcTkwV0jLwfWWth82pBceALEr5iCjY1GtYvpkxsOxeGEeEtr769ROXxO/bqfO1H
YfG0TU1EWVL77AoOv8+DNkbnYMaa53KjntlkrS4ifjZTVqLflp1zXTZwx7qBc0MlacIvgHMf92m8
LDKFvwunnPLryBzC6RgpLRbmZCaktkbmnEvm+eKWKstwru5LXyT9gx/P5zXzGNAJI+DCSXrQSYIC
Hd3Xstq8nRn7zdewA7YUBvEjCI5lb/doDZ3ZU9mMuQ+/gr6CmIJYq7mg9qA1etI4NOrcxjwcUsaN
ihPwou+u3A3c4ZazxMiK2I9MHbYIxVUblnxP7tIuFSkpbziiwn/aCVOHH6kNCN4W+TCct3YxiWxb
QUh/AhY1AA2A0HK7oKfx1ac8LuZiY3hn32KxspBAoIhMwPJ1IiTXV7sQaBVAFO5KyeiMy5n7jfb0
e6fDKeLgmJdUZjeUjMW+Y9S/s/yEuKVet0cYwHNmoBz9ChceqE8KJrS2opdhEZZw6s4tlhTwpJl0
3fhaewnRF1k+BBAwZIpYZfOhIwYrZCZF6Hnr+/NpVqz0oMwBl5WMKy9xznKZdS/tMgulDNTCBenG
vk5SwXNWxEYKfnmDHUlOwowKqKKXQRcJBGvDV6j1eh7/1srVZ2tmTj7TYBMMVDbU6x5veGGdXba/
QCzssR9AfmgFX3BgxcqrW1gXvA7t6beXJ6dAVJw3IfWZzE/JZM5KMuBoK190Z9TaUXrRFQv97k6x
C+qJqWXibdkptcrdV8kq1zHhWMrxLaYdY088Wxzwl8E1VwfZ85/7xIAN7qnao7ZNNW+USYN0fkM/
DD8vWBEifmiYQ8EeEjqfhbiDBtipOY+t7BNiXa5SpR5PEaFzEthGOswinnOLygBQXj4mrcbFhKi4
EotBqELQyVLgh1GVei5DQk85klfh1yprrErqRxx2kutut85H19bC6oOnVEEamJk697rvj1tmvr/g
DNnVEIi4JnoRhTlnXBjfz1LMspz4GEhhpYhHibYVJmKldDOr/5/QSSAtvTx6ZL4mwoPFZVTR6Rwj
HVxm/fH+DDzA/xDS0VPKNWH+RPbdzaCI4zlnyMsUit9tazs8FtNbDVeF8oReGKB6W0A0FSfQZem1
uO4RfFFoE8g1BDD+WPXU0k8XcrwYvo1NUw+3hDiw2m5Rx/rRv6x2IL02WbGI8UMdUYVcHwF0vudY
ur0q0FgnE1FtcK3OoFWHMiEHc19l8wppdXDifVmroJcvysGft62wluAtLm9ujk9eyhfixqCq2QZI
LX5EZLPt1uqJD6xsGO9n7Oby6ILxxBHX+P4OVO/+BzqMFbo2yMW/uOPL92I3Vyj6NW58vvYVJ+/4
Gg3z8xTKxDY5PnvkKGJ5h7THNmB9u+nyx2VZ2XyJnp7t3zbkg8bECkOQ+LfRDPJyfCK/IPxbIBhc
tKh88J/zz0sMVMjUjXlmGBxuexul5VMlcMEFYpT+hWgJi0XmD+JzyLykp94YOL2uSBYudBKTyqRf
UGgebeJbBevEi3bkUxvqQ6mmLC3b5MV9oRTp9dN28sqSUNvpDMwnF2V08XGerOQf5R6Cd9rtkbQ4
QMwAGyeWkkTQ0Us57VYFKNAMAd1ees+FfZedkwsTKYO/FLTojHxSSYjn03IeTmK+ElFLXiAa8yah
yg6EH5jyW8NsN/Y2U+AnCdwnXbxoZnb4vYHJxqoyLHmc0MKqCAQYzhX7Pi+1fXFdtcVYl/U7iEYD
Ht6oNMRX5CryDdzEAgErQVxSXSMyNQ2tlR8KgG6/zcdaXdk+5CYQ9ryvlolYHT1DWX7I7mj+fjlk
4oi1iy6t1g0EMwRExLnTdrZDO9a+Wa2cz8yLRC5YwMM//vmQqFdFsIEn4NunAWKyS6DYbYzOGm2F
+wV1aDqsaMheF6LJ6FEjDChW+Wp3yQ99VzXFHfctGGN09bi/Rc7g0HbRIU2uM0HK4uFEzzM72bu/
P93IRsm8cMkMy8PkRJuuuPPvnWzskLPr21eLdivwBHnjJwoG4pIbFWci8h1TK2r0Mpj7gh7DCQ55
VcImOYiO3ESy90oNVZpLiwqjXbOXFUk5Tj0Ru0g38PD0xvjI5vCxHJ3/QFxww2ID1jd7SoDrCUXP
d67Qr69Qmjft4y2+I7+zNfqWWkRvgeF+8ZAbbNFbmcsxoeEwxIw+larbwuT2KHa5zS2Jd/wc1Vfv
+ksJwW4/t5LxfO4i1c36YhP3AKJLkaS8oKcULUzyZVkmrEQ75f2pnC7Ee2urpSPACTEbbrZYf/gl
hIUu2r50ZgdFRLShI/kdPyxnO8a2rO+WAqTIe34kjZu+5QSWfil3Y2P+WgNUly2+f39RWvnu3y/W
5Np181btZ4caOjRu2wX0apPBcyrFSe+Bm0SEqy4niPomolDIZcjrjm33TFKfgTcyMyBvMxZjj0Jf
JwD9xpYTYSSMxrLrp1AGrGgKAElhZPKKyPtVlrErpLhBNrmTGu5yrp8VC5MB0pMXyFX/+5zJDyAa
3drseOQcp6dnHY8o0lq0OvR5bj5hVmbYnTVyBkiYbep6C6rDuksolOgdtJ3arEAtBF1NAeYv7CvJ
/2VCm1TqjGJx8oZ0NasWAXb2adlb+vgVp56NvPDPMGTNVw16ZVMq93x8jcmURexszUHchnkuKezE
XV0rISOucJo522dL2e8sq3GBKHO74SDf80pPS0AHAzyk9Hp/4cuBZhFe+xjFJm5TDATh8J2TmTvt
GJAuU3Nz3zEH97an3E42gLT/0kM8U9PUDY2z1wbGkFu1kDwcoM4SCp+c6wG3ETWHgI0ptXOnqPK6
dRafsTae6n1f+9TGop5BtwVm0sBjuRQdOwHa2mU0cccUQTMI31d8k1Hx6AYa792XdOBE05rJLufb
HYpQjbGDQlJOu/rRBUTe+lDOBuHbswXqE6OvfR20F1OxVdXzcnpp4JZ72/djbXeyIouVh97eWCuw
A4QvA8ME110ViCkMMDwoo1LFTzjjnRe+yGn9eoMCV2AGV5pcysWGLZUoFRvsNCWQGSYoNOMcRnai
KDpxIuQh8IYYcSgbki8CjPz4gkAmKW7xUx40N+i6k6m46hFQDCNXrjOGy7IqJkbax3NriX16nMB/
i7b19t5VsNKll6VVkoqyfCw0IuH4OSmW7o18GQk0By6gZTZhGGQyvI6Zs/tkOKHtJXS5gX8riT8V
D4QhaD7t4Neuy2Vlubh6CpeSP+p0XrbArWbPK5lW8Mgy0ZRXhl7zfTEGOk4Hwh2YUYKVMS/ijSDM
Sebg4Ts0lWUnmuMbIvkAZLijfMC2jOA4aXkUMZqNzU9le0mV3FsN0IAyaKmzu46Q0rd13720mBNi
EbAHM17h8sG4pI7dpMw/L2vcELxZzHQRMfzoU9J7snfusho3UV4BtG/jOFtxRVQvevVO6eLM1PXU
qzArIlSGJ4jKt0gEQr1lwNfqp9ivFFUWVE3OjJ4763XS+5ERTSbEUHvk6WFMDrfrF1BigSkenJsP
QDnSyvRXYX7g2rhNCfwRLE9K992s4FQ97s2WOnNgr2xtgn+e7JDzZYsiU1uNRc7s3LRJVSQLbpow
DnfEqlMiCx2+Ax7PQA45BX/qXSFsXjtNR0akLV4dI3XOxeUL08VM+ThSVXZFBDLNxsbG35Bw7rlH
SOGmHqXHE8H92Vi1Y4ypFAHXPp7oLFE5kqfxAA6DMEM7+45Rzxy/bd9xBoOQGx0b5qsFBJ+/VDw/
NYLweLykC8H/DtGFJcW4IMaMMrEvGoLeheSIaQJ12FQnsEJYaOCBDe6Ol7gHvBsQy6hT0Kle4iqC
/xww0AjZwxHog+ZroAi0eolPhvDj2Gua3hywCWLyyZSZzZAc85LtKsjU0/agrwi1fYc4L8F4OTcS
2Yu0JKErkJp2W7xBSPHXZAO8BX9VkM4ZTHxMRe3rBOKiHuLoJSF9DxC7BozATs4IOsZ9Y/14G/Wa
+/9t0kBbpSDWBnFCEyAuo5m2uVcyypzD0e7Not1Wrs+S4D/5e9qdq5ca+ITLcT3LE8H3u55XQ3bK
stguumHjuOvfwEVbC43f+Os0LXXkgWRd7N7hAvKrx9z+9enrG3MTe5OwT4WgL7875ZAMylrUiFat
viNhIQEz3Ie+Pc7tnIONY+jPgKYY8PlLff23S7PO5D0k4YFPnX/z/3EJ1omPEtrMHGx7Q176jG0G
JwmK+jpsdJFPhf8ygRv9aJ2+cBN8ku7R69mNWSUSksFqcjbBaImx84CzrIUH/VWtjqv/NSbLejgP
Wq3OIr5MLFqr/GcpJhSFGrrKNCGG1op+aIx/N2PQdhqhslzIw6ORtAqh0WYCV9Fcxekhhji9q2Ft
FCvz5eQEeXeSfTRWpG9XRy7fAGP0eRBe1ywFXanw4dinBRHueopukeHE9I1AqnmEqLHRwHOT29UW
CyEWjToIzhMfqovXFONEJVCMLwDwRAiHpUc5w1i85yzHryvuXbpEx8VA8BUMpQz+xPiVLmbmxOam
3Av3SB+FKbez1+5138/MCpqU336vpEEsszwc+5j+7DWfI5/PzFpc1LX1UOM64Cc6n6t9lBBeORJa
35Nx7xzcPYy+bS/wINeSyxGQ2DUjtyhE16x00EZm1kmwqvLtkPlKD4seqNG3ql3DbmTy57G99PS2
YTsb03OU2ZIAPbUnl+dAW5aZrgl9r57fFGDiRtZi7SwlPlaSmTmlGCQg+XEJ9xYbz3i8Q6+Cc1mQ
a+yKmp5jxamOkA/27uu3imWincXPtfnlKIFfVaTI8KjjXPWk7Wk8SVJr25VzVTg5Z9TiUIPTADgB
2eZr2R8iaAFXOCM5TndDE7MrJRHnybkWKVmRT10bEq58wqjTUAKmXd9gDrmF8YK/MkY3Cj+stfD7
2AevMLduQAhNprUFFW4BxP+ep1iR6KqrtredphKH/TYGHTjds/Mie1m3NiFPlxjpNFA62G5sf6LE
AM1fJVQ8nR4GxF/XRVaPY6jcvXQ/Hk9nOzziKb5bxoSdz2t5ud6r1eOz33xddCHWv1FbBJ2socsy
++os/aDYjJnUaAqZXB5JyXO2FADOcuUQSh0HcT5/NGL2MPIcf1wtL27M/LVssAnstw7NBCZWkwto
alHbJgeQHAHhEBFkQt9W/DvtV1DL69/fYSYqWKx0U7f5Fj2BA+FZf1PgnSSH6znj/e+RLZnyW8m1
Fqz2OiF9YSk1R1SDalc93a4471QrMM1G7toF3VEIMcMe/rBBSBcxTSCxNB83UylfMk7+YlhFf90S
iovi+cStLs6Cb60K0TTKJwGMo4nNudlAFETCQHETpiRKEwuRiz2d4zew8SgpBChXzcRvueqc9CO9
7ouk5rEd6PQqQjzbzHFfo41CxsLGnJG/qoiE3catIc4DplAHThhZKu+SKdDDP0rNGn1xgV1CdQZV
eEEP+3R+4G7vwwzm+vIXG7hr7lZifjKXi461sDUrClsKZCzLJTo5D6c7Bl9gOo6pRwh9nygSNbju
TYyWPFlBxEN1Ys6nsiAnViC0zPYhffW5WFzDryXKPKquRiGKDGOIfgxPBZeGjbRGToxyIUUn7haK
o6t4i7/aPaVRg3+e1iRnFRYgODPYmY7FrXSutbjzBsUbHW9wqF8d2F7S8MC1SJDpVBo5UveXYSqv
wDhfrEQXu/69qtteuv9mwRiME64szF8LR5fAlSmSZX1zv9vIxcZE1AVAjAk1BBZcbzMUboSdZWP/
TO/7aChURfw2dli21wFjZXIbxoYO9ub+I6EpcxQiSRTEtT9l8Xf5KD/GLUKl8ptDJOBBdmavD44w
N/Ipf2YN+yPjxx7gK+mu6Y3P33uGIDm1CswUkWkIOouIe4sj7WnBeyzMwyGFvB7JwL8k4H8kkiOq
JcAVFLIStKSN2bwdFwHnbt0fRibetlEmSZ+wMaRuZG0TnXFk8P/uBAT8S0JyvTpLM1TOpJRRd1Qj
tP+Cojg6qgNh796RswXy8tksWypM3KIeSCxg3X/qNC7wdeZRERlrU6cV1TxULzgTBI3clVW+EhNy
ehc0NpDzYycTRDMt50489Qh/pAFDtVcyRdIV9cbD5imxj6xRyOHkEHNmVsB/Ugt127Ae65HI3bL2
ePqJENuyE9BXJGYqURzn6RpyvxtIEVgKBnx4dFH686Bq+L4FfZok1GcthRK8nfW8J4TWj43rem9H
KPxDcjZnxO0+P3aGsIH8Gq1YWZEjcPdM59+plSkWZfZhggIXJSYxhODm3dbgSkgq6Dl5Bc8Qvk0u
RoWWVr6u/3rhxfIXo1ZXHselFem6dXKF2kjHOqxR1F2MM0SfpK/pxuW1bpKe80BelnQSYiAkOiCV
GOvynyh3Gwjnd5tNth4gZAMP0j8bs4BMFfe7H8RJQsuVEf4/vMmmxA2IgP5mj0Ag4XbFCtzFPJGR
DjImQ/pfaZaPDHiYcYjdBVNsbak/3HW06qbZiV3t04WKSGgiK7H88/p72RaALRsWfHkRhTMEoWDi
NFMZFLpqobsMMJ5IuYeRvL2wHs2RV6LIwSV4ceqt67KhIvilSF1wqFr1cu9p/iONi8s+ug1VZuuq
uPkPojJ03GIH6oTiqTK5krNu8xZNpzIgF98EgGjhesU2HY3GoqfO7j6K2kU430LNs1SLQS4DIpj2
tSGZchMBz07K4QoGIGsmfDz5moiE02N9ZeFlAJgHDoRgNzDpB0ls2q0STLdyaekS0d0BrKOmEk5B
eVBZDVFVyux3DAX1PB5QZmnR6CieFiFUtTXWyktxYUYfbTy7S+LuAu0giWX2iJ//nKk64A7WyRVF
uMjVCS5es+AAKq/24HFqpoUXjx3rAaaFKDjbmm/eyz5fUcv8/XB5W26E1fh5Gc9E1j1gypQ5y1Dh
y53hCQuPK5nsYv3XtYSpTS3xddOJl0CNtJOzUTToZ97ww9jG5xhjmJ63Vf9JZXXb+f/NUnJVGqdQ
nBBhz5iZJCBGopl1e5yjYWXj1IbvwXk3Pyr4+k/DtrnghrMvan62hNqsvpGpM2KAefW1pVPVTHKb
g0Ut0upuoLM/UT6rQe791y3bJyoxgiWOeByJ5cTamriXRrySpTFnj7XimPsHv1wVDNo2i4t118ao
KTN8rUSrQXRHQOlMn9g3sQUy18MBX4AJg+aZ8VMSGMX2bhpff1bS91EF4SzlP56D5Dhp8ArR/8Ud
w6VZ7Zq/WuOea/9xdd9kOokVlljrHkwQjG3PVR2VO6aiojRXv+uPy19HUsaOq28mAmH4vddegfy9
eW/Zp9YBIIHEkat6TH1ssLSaQoShoJfHf3/vOLG1R60vcAiXsb+VVN5x6M6O9HsHXyO8mDDh82wQ
bCzWwizk7QqpFqOdfl52dTqpHyHM4DgKg1cEJ064EcOZ6U5D/DpAlHX9la+eUhesFvhcMu1jkroD
LGkpbWMdu2Rw0Z41AD60sXHsv45GN7oA8FdSipiL9Tqs0UB+S+1iGYOBN9qS5SuG19k3cBH4FZ40
K6+R+4uR/RnUXNYAvFlIeWcbe8qGWQx4E7SDdaGFycKWPgIKzWNDuJjK6UxUOmhHGHyqrvdX8kUY
SX/eFSIl4AuGkZzVaffYyVNFKmkWXsqjcYC93zAEA+o8V2EtVB1ADvnBjjDkzl+l2CUmQFODv9DR
Yml0Yw5gWBvcQXkuuAnBOAeyieJHPMXnFVxA3HZldHy20OrTOsUXKmkSmY3CaSkg4R+QD8scdRcA
/xApx9Wq+sFzFeYg6rvvSTJJfd0ZjRWhZl6FJdVabOM1C1ODtut+XQLgREUPk6QtX7eEbObTvPUf
wLffgKKX2YbHpoYlqr3jZh/nfKtCNxhpWxLtwOOUDgua7IfCQlCBrzDAi2eT4btSh5mU8eEV33NP
3D6X10GOin3gWr7V1byMCofqV52MX+ygy76uRvBrD4M3boPOfH6BJhR+N1BLb8jSRqQweI0JnxAN
QUtq9fIz3ZGkYVrXjxmG6Mbe1+543lU4tGuEvvHVzK/nscqghyJzwARh+xQsq2Rl0YXsW1foNMsI
0Q0PtLH7vHMfW/ZwXzRe7shNSyacGliQEsSfGdjheYkRagH++CuJEKIRdHez9tiDeTh6XqGVoJ+F
QpnlnXfIK9ajoJnUxHpoKHipEkvRZnqJzU0GqOe01NJmu+7trIhUl3u9CQX6R+o/8at9B/T70SCm
qFScR3ePDS+7nTQlJ2kBC3rn3zEQjcDnSu6aNjosnOcFYT6uNOoMuTRdqzZ+KEhjSVYEnKKiCgPo
bWqm8NkyXepHSAIEswAY0VIrl4MURiBw63m+6MB57TiBKZupu/PHn0siYKiqKZ8VcCQAg4AfCGUv
aW+R8+yG8YgHXDCqoxYi3weapEqUYn8fm/6DyKzLqbxmuupxa1bTwJBznJadloyDWVjYQ4cg3u1o
NqyhUV4+maxW3RfPLUj6grgm1jtQfJ4Cvno9nkWIvdPc7icHI9ktkuwPWLNdHiL/uhRGzkP2qI2E
iamHFCnh87psM6OSJ41TflA4YyArhJNN3BUEZVZ9+vooRzzWosMGUP+7wTpkEs0WisyvnLiihHPK
ziUhpsEQUy7K+bJlA2HVYiUsG6oKXZQjdB+vtmSLhkz93RZA0Oqr5lKxx5uU+/ljAd62lyH7gH+Z
Qkrc8VMjnqAdiQUWeHvucFJb+tVbVG1vivW47vLgsF8rzbKp+ztGZiFmRqTysHkx8xdDNvkpAu6v
XAweVsvpE/6SFyDz2w3CyjL+Td+i1yOn7wKvu2WCaT1HyLwSqMbq4o9uL7TpqaeOTqXpESf5xAQo
SQqq63fFzS5P9zU1FbpvGzt26hTh4F5TQ9c/irooDnlOYVJC5Q9bHS6YpoP/rMxXxPj64CY2ntNr
NHGgzUw2aZRob0fGHrSrSTHjiY2KJ6zsRlM6MgD1kCGOkiXczB4xlD4+pXuF4sWkRYg7Z2MYOJcM
Scwh2qcfNe6uyxLKq++VnpSNyDHHe5lc0o1ojrtTi/5snz0aUWrbTUxkdRCz8UJ4GDhZ0R5cKM95
2B8qyWqvwqTuy/Jjh+lPboxwWftV107tPaN2JwtJREvWG+vzvtS4pdIPv0+KYzecILfDnLId2C9t
svm8NA8/5bM2nsaOQeRAZkLolzDiw51XihXoW3fCPz/pYzeaSDfiLtCGX7iSVdYDmOrOKfQ/CwTI
aZkhGfu/gNJiNPJR4gkYsBVMJSfYk6Qm6mthKrwm2c52fYL08FUlyttAto5fKWNgicG2VVOvZcQi
8dqYZHuXkS72WCj0AmAfyxDCxAWeIe2b0S/Rc4Gk1ML6/pnj7SwkD2WngC5+JqoedaGDT6UTE3Ca
lfkTSOPHYcU6XvgrC6ofVKs5LByxdNScFmX1df/ZVrxEO6HG6isu+iQwjUmvHLkMxjslKR4qj20Y
/dnQb345Jj/EJGCUJGIiLojhphk8Pqtb1sMZYYVzo2Rftu5uBcF4RKt/GDY35Df1yYuqOcS7lxGJ
T5lQjaSyBBSusZZ1Y4y6DDSpGB1S2o+PRj1q4XZZvZQ16KgvqbQpq9hxUjmRNQaiomUIitq/M/xS
3InG3R8nfCJwWeeKivhwcIyPSr4Yd75gGwRWoZ8Sy7TKCVo9j4vKIwIC1YhbArkTU6Z7uwhw54Lr
OcoivQwVaTMEzo53VfS2lvjYHwI5YBO3aF6TUBRG0ip4W3z/YXeiGT2D7MFW1fkELAytK8DBI4my
1xxIIgJP+VRi+bRt9oWtm7xL9jWSF7EbZqwsfcQ8zKumEV8CWctQ2kVFYkhb5wY+InN9xOd3XTL8
vPE+MearurxaLYPqHBkTRm2tBo17uiDqvnBfQKcfN2afOZ+vU7pQiVhpotlmtDb/HjaoyLZekRRJ
7YHS1yaeklBTaamLF4AZ9YFf7m+3imNQhAmlzErL0cJivAEBOoEUBsN08sQpUyVCqTamcWWC2/md
dd8QxjIbtBsUNhCqVJ4t026O88piKl8mz6VPRMhNdZk/3BzteregpCNXm8oCHAJyUmy4Lr5Dspe6
vL5ob7sHGwWkct4dU6cVTXQXzmD4yrdMvVklmChnYCaHF8O+sWEp2s3yaJvNwOYvE/gq9g7nvYkJ
+CoI7Uxnlzsx1dmqZCVlakykenzHqWj/N8MGdpSka4jadpDen7DLgqrRNkKuw7T8i29qwlD65iqH
QOCToyBQ8b/kbPezszBS2j3VMYTurfOsu2pxT/FqZwjQYUtxoBwdMlisSwj+debnyfUMF5F3DSY3
29paeVHOyVPX8UiCB5JvlmNmuHxYb+3K6pFiUYFk6TZgjYsgG8Ex8qA7hq8vLFEkGzVb8+li6+Dy
DZeaY42XrRGtdns7hSaRdX6eWOF6jYlLdzDUmNEef4MGPv737WEuhwOOwWTG2/dLVE+ZLDqz1yp3
oMVOdqHhzXhxRCEtsnoh2Mii3jBs+9Vi7FgUCby/IQDWFSuT8n9k6onQ0UzWOSAQQxXa8F4mSbWd
yHuc4G7A+W9YnGFAval1ZOSOXoTW24wAUeJrsoFcuvOMzrKK6HIt/bzyEQ968KwnldQrclPQcIkr
nWPWSJNtpCWWZqhUeSDGG83RJoITtEb8F+HGWqUpGSaUVsmfc+tf4MRYTSTAikngwIFNdrOkfJRa
2PJrtNcFvMOvGyIq6DPS4Djxy0oylof69yInu0tZzBbCZBUcGqDp1xEcGezbRDks7/AzR/9nUt3G
FJ3E2267jFhYIV5cP1oJznX7AA+TFIq3FUHCkEwZR9xQUMjbINk1+srxPa6T3/twg8EA3NrQGZ3e
x7tr7naCuSxYQbipxZdE/8maTYoWRdCK5j7saX3F4694aqpY13XgreXtTJrYQXAcZqqQH1xkhI+E
RXDrG4cHcT4tN3BXKQ3EUH21lknsFBI7pftjOva36Dh9HRTM6oTeMJwoW+C9Pm+PhCqSv7HMRjgl
Es+fkR6qQkfbpnD4XZ9kMWoEJhWJR3ZDI4bMWBf1Wkqx4w5xer15umDXA2zFRJguC7pKSnHdVeaf
VVn5IwJgsc9kLRO+1QCRxUPA8Kxzqd0iEKpMdinMPpWMpRQXgo+mu19YAiZKEEcPpSwExQAIxdXC
ZEIKultDcIw2pFTYQ6TtHVL5jW2Obf3tIg2CZRnJyzNbxhePzmHXjE3RCtR1t7AgzIVzIEvHdt90
SL9/xNh6sQmtu4fvPdAYTzGCAF5Xn7/NWp4UeIirtvd7OkH/R5VKzsF487sEXzD3vCc+mjqqeEKL
3mKBtrQqFLPJli8GXManl7zM2IBbv0zrEgDMzsKwhuSgg/V/FFwf21yO9S2PIquQDGg2wg6bjver
4rEJZ+k0osAl2hqPB3lUaVwgm+O/bQXiqtIaLWQpLJVoWwfSxcLnAQrqP6uTY/LdquViexlQw6vN
AXiyHHDhZsYHRPHrEFXNGsL4+6ppvvqTMKd/myUf5Pm+s+VrqqDAG+pspnnaK6USWGo6HjicvJ4K
GYuxLpY7IShAKxW0f+YshdCJxAuxueJs0hIPcfWp3pBmQc/RxKXfjaSN1H72ykN5AlHDRzjU+wYQ
+/YSTgFC2RT3S5XYSBkpCDozIbzv+hrUwbtMkw3r9P8b9cfNFNKJzqi9ovnCF1sCuXA5KmA4Pvfz
V6LB1UBkJd6cDhUvZeoRDbjaXn/f5WxtkfVu45EDWiyaQHgVfF+6Ra3YDm719Es524Lt4633p9WV
Koae/cJOFru4U9FTfb6X1CyNkarZBQgFDXRW9/RFkJuNibBiG/B2ORbB8jg5dHoVjH+wivwfa7vZ
ucaxuBeATlxJw8BepRd/JeoZYBugQXTunQD3qIYW5RHakl4mIqr6bQD9KmiFGfR33+vR0rMAWjkY
1AeIxf0eOjOJRA/Ga6sQX70GWz6lnzX96wiQ4KtsYJ9RHPQyY6EAWpbj3LtBG6LUHAmS/bvTxWi7
/B4UEjHXJ9CuINqDQc4W9F7CbZhye/He8wrw2L6a9QqKe1bs6uUJGUPzq8rGIJA3CCNaxLiSOyUL
rUjLlesBvZ/1v7xmrzo3WgkLTWwQlQjB+qOTVno9cp+q+j60WhZ2y7ER5KW5wgvMphZ4AWTNoP3o
+5GpoclxCiHftqscISPlnKkhaXZxxg/SER2vMwbayfiLW+W/q23Ovx0waZwe2C1VuzNCEV1ah7+w
XcG10XHYbQJMPyeAx/ek7XMdgfJmocT4OQ+OXjqqjNKX2syrja8ic39uf/9y18M3HjShm2GQnIZf
DfXinf+KlJWwXYzC1ZsCNg/46XEJEdYhbAG1U8CHmas1xufeTcOq2/YJcTbnyGacmJliL7WFhYBq
WfxJTZZ5m1AqPPURGiMKThAIn4itxDM5rsc++Y8o9FMJnCj/CU8UUxPuwgkOAqA6ivB9hJ9SOHrn
st6Nxbtfbwh7YZSpe6YFUbh/o6pnVdS6SB/KMD2NnsvxyNJyhV8KJtE6olXUQVI4jZtGI+PqqP85
vj2krWwvQeEC/SdjleLA7apxxBBDrDGZSfIis12t4KiLAVOUFqkq15Et+g8Cq+jyylZKgz571t7d
zk5awFh+KcsEPaudImBGOAYoASPtWIMjWRWbGHC0xRVOrQMZoB1R3FY9sAwtVhDSC8v8sacK53ax
bGkaoP66zeIXbubxna0PZrZm0e9txIS2T+UxF9xtgp6+2lipaMgWf5LzEdmsfUY9usrbcsektUps
m812ovF1QUxU237P55Vv4FcOltHI153h4HMT/xLe4xynqK3Bb8GRg9XSTui92HUG9UEoMioJj1hE
ipT/o3ovqitPjq6t92kfelaCtxynUX2ncAmDIpG/qDGNTdNlzkX/x35DPvBlqucPfARGU5PfDtVg
ELFP+qwzvnXL/WLuRj4MILqaq4RISc/Ew9rdaSrhej6ilthLiMW1+lrnKlWOerUR9JqZPI2OQWYe
jUNJS1LdJBwYfo6rK5vSJJoryiSMyV0m3MMUMuux55G1ROS8tDQCchiVorf8/Hw93XVsOLtFYBrG
qmSg0ZHbrcsH1N/Mdx9ioZn+73mDQGdJzEpdWJwZbNc5ZxE0ImilBXVg/qaDbCRzjaDAz/SEGHIb
W9MVOLPxVYRuUs/F3sRlO20fa7YXmZlknAyuXGA07pR9G3QHtmLjZ+8YacjV9C8QgDrGs5vtwy5e
SJGfwm3r3fTEdU7eNxwtuY0MQmPNPaC2dcisy6v29Iu376wes6EV5qafAwbnwq8EV625X0n3s4ZF
Zt95rrP1vvUWvoN24UEBrmNCc75p0nS0928QhMD4PmO8Isrn3JHS7FxmXMLU+ba3nMGVppxwn9+l
jmeD5ZU2jmPXIis6bnYVs0x4V2CLnasOP8JoNi1+LbZ+hgHEiLZ934KiXWPRSN/Zd46F5gPKGmRh
GjlYdleNQOoeBbOuyHMTKsXBOWMZtAskz5Wl2yobWnpbRVzvRBr3atD6a8X7nDQlA69A1OVSCbYx
Mwosw17rzzU2bddmhrwQEvPOC+jQqu7WuohC4uabe9r20UCq1wl2rtnLw9VODUdt+wPCcivHSRBc
piS8YTuht8/sSrdZIC2j6cPSgwe1tesx9laVy8w14+X+wsZhyyw68wdDP/hrVcBYopH+jbpMqO43
sD3VimuyV+3V5U0A31bNzd08htK0dhw2JLNmn85diwMFTZe+HiJB1lVjvzVaAAFTRi9Hqku8HgzG
ayaKy2sZyWfkXCfB7fapgOE4m9ddA63LudhRxnTw7Ej+vK9z80XP1r1HYUnXDCPZB5b3t1rNiKLL
1hvzDM2jvicx0mN/Bo8+7Rt23ARmIDgDssU9Hby6bzXOTUVZUCjS4exRUQtd7WhcYgSV8721DCxn
lhXVxeTtbyGy2c4SYg9PSZyt1flmbJ3BGqAdtQN2fO+qHAhgOGfCEU3l4h9JliMXseFpeH4ompbk
WLM5x0Cswv7FRstbcnpw2roaDhngYLVbjEzbZXqlMSMw6LxyKEgUnLcc3adQ8Yw0acspsrkEyP4l
FQ5dXARr1F+69FhjvQv5aGkD864iNr1+WUxYBhjpOdDHAGRxQXvn9WFDk8ZHwxxoahtAu/Xk3JdG
GM53LKL+8D7mLfbW2E/CLKSp2EJI8MjHHWfX5w+KPPIaBs0JYNY6yF1fKEDm3FoZ0efo9ftxxaHI
IcRs2j1+O0hbtYEzP4rfsvgmEgdriuekrevZF+Z9TrB0n5LFQgSaZIa8TONV4Tb2wiV4wTHGOUW5
aLfuWg2hvkP7gUAZHvMz93RkEso+2GVV+EfNMgG3N4LBu20NswrjT6MXFpOHKGW/+ziQ6l3dQxK4
ElbSK9wgommLZ4ZABwL/whj50l+1+js5g5LwXcp3YUIUJvZkaLfoRiEAMOfHrE6p/qtwlL71nXD3
48T4GhAq7iIUOwTiI3idsjB3pUBeGqd58wsNDRDTwFIbK1bJDhUQt+ByCzszERw78Wdhx14QArwK
aEyEexLxnOazZkCHuYQDsXOkJvLSkIcEZhHjwE1z3BsTbDg47TbmtqZ4xRD34As8YPXKcRqf21lY
/fs0N9S5MTfd2Z6Ie2KOZ5MKSMspXB7w6M6MddtSt/UkzDIFmQC86g6ADpQEI+Jl3ertIq0focwK
G4ef8QzAAZsWxr3YhAQJH7/5CYkGdVGXfeU/XSULUdIuV3l/NIiO+mgooQoEcBMLR1akaytRajVy
MGG4iOhhuqJCasDrHnLmdbiGwtHRgPe/TpRHuFNs5bFP5T8M4FDs7oZ6IMJmUcdyGYrDbZ+k2EWL
mW2mxMwsZUCnkSRnAO+6caPXLEwwrToPsexmJioX+m+gHLhIFWkkildEVEz2YHlCL6Q751K/H0Iw
YCwNLrEVDdj7rjm8/jCtUxxSCnXbjPEO+zi/YTwNliYJFdY+ZvULcgkE5eaa1vXlb+0VX46P8mEn
ODgGsgoh903zfpiay6Ua8v7ZQ+q/ggqyRVZBTXSQ4qR6XyB6zeLtUYA6h7OzvuvBxAFLYvBGd7QW
cQCPzUDecLx6Onw/4S/QC4Ll3jEALDk72LDhmNLZsGN4rqUGX6pAGc9xbU9JKjfS2p+AgusEY/79
uSU/qSLuONP4hlurT80Pk2lRbQskh2VFSV9xHQtuVP65OvqwPb01JmXlaYOUe029G9XwNhXx+ma4
ZyB7J67TI+4ebVz5CIi8DWU2aUeW9iMpgVpm51jxT7XgHhkuukZCgjcVDlg7eU/7UVsapJxDOTjH
aUByM9NWx2k1p4qszNzV4RqmUsjM6bwxtx+2Rd9oR9EVshrXWXFMEKl/OMD3wHONVCy/qIrTBkWa
9uhGwndHEzIVgg9rPD1IZRIavCoGGohCR7JUDpOIvlI+i1rrDjbpJWcDYuFoOkynQxVlkDRGjd57
NJyNRmZZCo8i4mqaj7p6Gv91rrNW7KbRB2ltn1VY+udPMrKxGUN/Q51I8eIlFyaNm9UFyMpC+wMJ
4wH2Je4EJboPgghxz/6JzJJuSyswdiGQEnvNX1TQKdunpjQQJ1zvzNY9GKhn4foKbdnVlvXqPcRz
KFZ374C+qfGJW6iH6xNGJnFgjTJvQexy3DTsG0kewJoBHzLsNODv4sfdq2tH4qQ9rzWvz2IJJwAM
xRRxZIHRibFyYGEDeelswW8xbBrRTtRKf7DvHgG+b23EBHCotDNlq5VtbdW5Vwa+/6PtGpJc5N/c
PufaCvewXz2fk45ARmJgfaUqT8nEaQtjzMaVFkbC/VIdtVtBrP2wasFtdL9tVbnD41u/4qJ2wxqs
wXlLSnWorzRvmezaYiWZlGdeCi13Kjhf9FeBEM0LNEMMpxbbiyzF77QYoyXAA3W+aXWf1Rp1FgsB
dwxB4gZGmE69KLMkK3I5Ntin/8CCVc2olHW30vjdK+xeEKer3NZDwgSBL/W6QYmxQSYHXi3jijAd
Y/kETj7baZ28pS+SIXjB9DHB2lB/GaZqpddGMcZHXUjE3yUnMzeVEyJh9cbMaaeZA+vo838nUxOk
XH2/B55LoF6bcQOS5ck3OAVYpcUXrEk9GtEIiF2bfX6oaclUvjJ0ij0UsMXv9eU2tC3T6Vpm47Ve
HtSh2grxqce0HJacDVRarzdlcjNv3eBSvSMg8Ir4Z4yIBPcAqr3/49Gsa1yVaws83M48aooIB90E
w4DU1cGJIcTelbycXJRj4RRccJxHDBI+ZmKKaHUFU+FiA5mL+SThxgp/lDA4pQw6a1q+hcK40wTw
IIBk1usX+DKRkj4mVXa9cO26nSuebDHzTEzTrkMyCge28AKbRe2AHJ2hxDJjRdQOYCNP1s9Z/Y+p
pS9S4pfMatTtCcZGdZqQPnv6w6WABz0XjEmVfDrkbwlT9cZAShAC8jDEkZjklrnIhvIK4IHTN/xC
wQtmt5S4VzCXSJEqZ2hLEwN31SmhqnOcpZrPY3aHATW+bmwzLh2LvSSu3NJ2YrUbVlDH73/FhuUf
aDOmBVZZ5g7+BTgWRSh2n6Tt7LpN66SR07OyAbVO4TuRw6/fnipWDF7r8mXsCnOU04oICw5c2WWa
VdTD95AXaad5ZXQ3euhElSlD2BxK3bPdOgqQYY8ErF7c80vr0Dr26nGP4Ruc/jYgaZh5NdWwh69O
4l6a/JRByOXGODNlZLehR0csFEKfIH/Ikbdi/r6slmgs+jPo+Ev5oVhVHhcELc2ZpKT6SPNtlq/r
2xr02TMv1fIkpRzNTI7nPN4KaZljs1+24HMXa6XFQwnXcAEXdnm/ZFFf/pVP4+dw9cYWvEsoEtN+
pIgK1WBoIlpT5WKEYdHq1qWsCSTeqB9fLFr3L6FmOyi8sgRsmAFoPlDxW6F2qAY98s9Dx/sw9t77
lUx3ymFmg6DS4dT8uakeut3LZZgcnuYEXi7X9fi/ky8LMyRexEFwEdsbLF094WPyu7me1gttRZ5k
XibojgjUOr6BZCbtma1rp0fKhcmjwikUbd+HFNY5/V1etbnsejnUfJmCL4VL1LpfpT+jx7baoduW
LMXqz4OhZviy/k4h+fyt5xmNopNjzgfrt+tnA8puzbE/Gxu9kPnnKymZYAXOLz0vIhFFqonVWXni
D/Uthn8HVm2w3wQsCzZ3RpkObI2D9swWXVFHk1EYCG255zZgBZ7XXx51HxcigO7TUUsmVgSH7dAD
1wYleguOiTw0x4gjSbp7BJeovDbcqPiTPTypagin6/sbd/8fxODhwh5f2tkO127GCgA7KsOG3cjj
XqDK4YQnaRCNoU+wrCkPyI9fykrDljCKG2p6cfMBGWorgP0zzZkiDzOgOk7VUphhAV5KoOHbOWAs
ANV4ws5dUDxWH3ZYyow2glrYMws5jLuCyo2bmlJkS5aPEhJVw1LN37FygcpipojU68lhc02mK/m6
GAfasb1WtgZk0J2idXed/c/JWsTTGBgkp7iZX5Qc3TK5BipbR9k08iqhyMSxH56DsVbSkFi8zNF0
O0C6vC9IvwWQSRtbD7B/ZSiWWwZNbg32amOkze6bCLYcfkuBv1M1x8px83mkMkSoVEgVQcWz8Ejd
3Iic4035K39Vl0kjLvX3iWnydhZa11KaGQ460bB8ardeyimKpCMq6s95sYPINf/4JSLOh+Ic/Cn7
l19DJSoRKDUy1Cy+Uwt0n4SfJErVZ7N1h4nplp69WrARBT2q6FPX1ljSiKIqmze5x14xdQv+Q6xU
97F/Kb0OqO4GTAYQfdH8AqxntwEj2ov3C6PgLXbVmpNvJ3MVx3RWU9lPpDQ6lApq9dmRDtfA5tTh
/6wE157cY7uePLaHFOYszR7g6o5dluT+6/reOQYzr/hPwXrnDIAZTx2gjLPIZv9AQRmPbZS1CsZN
DO8hJ8lrjcz1doMCjWMjrRDKpMYaD97umWW7WsmI6jv6FxDhYe+dr4ZT9SsU0xLWOKycC5WLfbDX
BYJQFH1dpLYKr5vSP4kYXY0nlIch0ujIAlL2dwmJnipIVJNQ9TLmh//a1jMoprU6j+IncZn1f5EI
uCsE0+JeBdtVZko7oq5ARp0EDP13cpQfv000ROLDph7KpecVKAn63vNQBQu/izPdVGth5jMEhCd9
QdODZFg8zi4XiMzeP3K3pAViXhshCi6xMyekl5Fpz0Wnqw00FGEgsz3pwac+vhjptsqYLv7nwIEC
GtNHVRJgEHdOO/FLvD0B8ka9LyNNccAEF1+pyVMIARt2myCzt6Xfb2dMniSgoZKMQeqJ43njQO5z
nCmUXuo4iCzHovMiK+tjLVnhCPePcfEkCgX+En/S4LbLqtabYNtqDWsY3qOS27GqnSr2Qw7cEhCz
hL+/LDeeTrqkjCHoorafyofDg1xLY464QzjMgqps8serVjyQu6wBoCyK6nzKmTiTcwwCTBGM0NKN
8lNG86JGSqE1zeSL6l6lQRGsKlhG+yif7nuRSW/et6IlfoG28fReDtdyTHQLCzET6b/4J8NK/M6g
x+r/pSLG/6VdnOwvKbxBoVvUYofftaS1gCoAT5vFCaxT7xL13YMdOkgBjZrmZn+NS6pMQAnK8xv5
5z5u3WVdksQgPlUQJ9m77NPm06lXUf9zmZmNwkPAfN5m5dk/4RYGExKUMlzyesjeFgIzs9unUVq/
JrtqeCwFWkWc1n0kn4bwEOqob2OCWHVynMpS5Ppj4QDZsT9eS+/ys+gGjsPp4iICvdBPBLDY1w5I
OtvFt4RRrDPZcd+10qcwvZ7TTz+jogmCyzxTBPZrgQA031LlXDsRpmUd0Gg+Vcfpe2zBBxzNAWnB
K91YvVT7UIrgRHFP//1KN6/tT+3fUf5ai8ra1iaE8gS3NiHjrazEzsaEVnG3Td7tYTGKdQKFVPaL
J/mc2E1x+LrnbkEMtL/qBczJK3D33FLIwROgMNvgMZ9sR3Js+BB+m2Ly7Iza+rsjDNmOFeDDt97s
Ajv/QidxT/qpmY/CLiRDfB/P+wStvy33a2tXb1mOq+V4ZF34jPvYNawWL4B1lyyzfQGZUcgXImW/
v4KPpQBNSBRAxgOKlSrR13GPauDPUfOehW4etqsSM1lNehZcBMefzTwCtoiTAwjiCDv9oAGnMhz4
RadO0DP8q+Nhc4eW42yERs+SBk6B42m8fKy1G7jkFG9dwcm1hkZrGSEckE8Oia1p5OQy7WLVxEzS
Gu/KJAkZcsIcp0uHxin+iKoYaJfB4Z6S6lV9RuPTA7CBdhlc1TX/FHGydC6QeEG+qapWiNPVuhrh
FYr52+sQ1Zv7gAnK+0yYFmvqPaNLWnxbV/Bu0T+99Z3cwGM7Jb4+UsbyoaY9C1jn1urvyhlKbuTB
pV/dJE4L+jzRxQHgr1ef7E+Eu6myl1pj+USAt1e4Ok+q4rLSjvkebib7droRY6/L2u9xHrIti53y
VeNrP5+9SMyQa2+ayHeXnE/dSrak94zE1fz2PM2x0utzGnvpFEkIipYKWer8jE9OWeOGDeZzATc9
7U4iVniMXBr216LYUrS31DSQhxgfmPiHED7VEce8FYAc9/hl6cgbwFacoWL3CBgqlaoad/bamser
Ms+rG19xgZO0LGjLCoZ9+SHbgFTSe977NIeMIPvR6rlTo4RG+SZMQDoDgoprguveqZmNql1QW7U3
A88wgFSBUKyloQWloZX1Z7hWEbXElVLkgvbK19mimtwKPJxci4RkmI9j9ZeqdgWxXgiqNER19O7v
HX27oE6x11ZFFGj6fHuor93wN2W+tcXBWqhUqHx1a4bNutNr1QnUgzRqhTX+q5AlkA3jcL4thso+
Pig+6WKVuhUNImEN5RYTlDh2aYacvy1uhub3t7jl4AIftiyEi2yHvE4OiUG1WLIhh7HUlnZ4/K7F
7Kax2GphvbSGwYXXcOGDEJX5FSTxP3tC24b10d3+7qAKdZo1xfsj5WftWaSd1pbgD+687L2q9dIj
rYlAb7CTEVp/XsqJ6V+RoKbGwreggDZ2eZFEoh0p6WvhcgQvj+i2ElXvBCVgur6tkMKNf7Jd2ORd
7Nm2VrC6o0Qdjhowzic7eW3zzSyyzgLs+46wSjHL+CDjTfd1jCYvUrhWU22wPQ17Iax+V7/Og3uF
QJdNmA3VhsEryBLVLEN2qTMZXaQvsvFvCza0lAMfAv3u3qSweL9sydC8H2764eFNSBYiggJLiQYg
HCafcvrC9mXV2IZGSYrPn7RWPF6DcJ3H2+g5G6+duhLJIi6L+/wHwp2+ndy/00v8ffa9ZssbUZO7
MB+CO22U4lMHQJl21zJOi7WzH2n6erf4Kq/eWvSlX10O2U7hldEwUOP3nIz6ac9aQD/bhAHzkhgn
Wdv1MpVa8i2Oxb8/nuqyKWMOdxtxyYsYD297PWsrIJMgcPQonQwtge1W/qtg/AEVtuqGhlc6Q7bC
JMMYqfBya0hAfSmnWSJQdy0py15NOEmi86CL6o10nvtl7z/lrQGY38/UpEO/buuO/hVXuYxuAef+
DADTBKTYRyNMdsgXF/YG/ch8Lc2YB/y+725l/BNLGQuw7Z8+5sisw6sG4woEv54auJR4ieGQBSR4
o9HpzQNSwA1ctV6ESY8Hut5ocH+Xx6h59rtAKS8DJwL9PewVUD4hq78KmJ1SrXADefChhjni1MpI
itzGMRDLz+KV1elpNg1SfWBeP0myeKF+1v+m4hmUq2j9V7XzQcQwTtE3++WYZcmZgCVcO3/TWhiA
LMV9sLklARWepICIA90MajEPK0peqG1K2S6DsBxvF0JI6RADAin7ROzLH2Gt0BUwG2vbeKM6jEQX
VvWFDHSpYLq2dzhAFmMB4s9+19cGU4LKA8NAOvwxz9f2PvBBHK+TiTZgHyEDtmK2X4a2SZOC8moX
wQa+EMf53yrMu+ESsaGlXZ586H/K1Q7si4tLnHXuvGjiqgQBzFtWMVMJ+U6eprxViUEsIqdUQ+ZH
7nHnPfjNmA2K82QsJMH0fanbZSIVsMO9KOL3oSHr/4VzVJE9DS4tH3LvtBuNkPcY92DlvFk9ozhQ
4fngAo4hzeb2M2RrR6W3C4Hfdy3TkOQVDx5YojkLoFBjriqLnnzcf5bgBoTqbWPMhSCMhkKhwR3d
Czp4v4aThv/e37/EnvuzoRAamTgs6BLPWsQ29WNt8bSFk6tFhF/ttUKAvERenmguMg44Kj9VoKMr
LCVHP1iDyllAAd806uzEQoxvEVVv2voTKSG3Dw8QTSxsPVCprnSy9EOSyo7Gj4Shcf7LsKbtYXIr
6Hik1Ea1yVoXi7IJcqf4xJMmdfJxsT3vC71oNjLvnuLI1iExRzLVTlnpftzvGPyyRMSYd/n2SgOX
MIEN1tPUmcyfxONuQR7VQ92Y5iCil1u/8dLAWR2v+bShnZhu6EHCDbNTIstHEt5kSsq/u4Jbj4RX
3VJItyFGyETGK+NxIYDmAQYEvGStRWLJoI0Q2P49jHlcG0AQHO4nj3X+r4RIA1nCFFuA8sIuD4TB
URdXBoIkLT3vw/CfBmAklc+8HqRRIN/nkwAXBT1akYwGHWELZaEo2fziwUNIYq3fm6Vb1ExmbFeQ
tdyoXjdbgHILf4/IUPLIz5NLWuyJeofBW0azdwnCHl9BJ7MpfLM2qP+86+VRIjW6ULO6/lKL+DYb
PFUmAe2jVuhoZ1aRpp+4YDTGSba/6KsN7Muae7gzM8k+xOwPiflg5BqHfUSlNJ3i7Okn6jn42YUk
ugjqdUOWTVDZDCWJik7ze/s2SbA2HmvyAZMCoH6hcZyRLjE7POtUWAxjB7cuSUp7zCu0CfSMRZ5s
4Y+atcwl67lJUG34aDHvoI0+tNJZphncOd5KW/kiS81VTleWBvryzb58wTnDJ+xpd4FZTvwEuLDj
1RsJOy4Q/cFAoyVS6UKoHtHVW4p+ZhRqx6ulr+iWY4U90iyR10EkZJSJbHXNROJzGx6pBcrUlblT
jIAEzBrDyqaRlHjfZJkqk95JPFwSGZM/SN7JHjYADNOR9mz3oMJHC5lzduL/B4Tj+eikTiBYrpB5
L8o4pQ9+rV3QGVeTA6Sa4eTIE1HephWuhMPkzYtVrpzgfNwXe/jpwvRYdsYPWTSEPuEEnI24b+eD
biTZGPhCzyIM2oteLv79aljIvUn3615nxjJkhbJjXCPMBGyLUkoozPNzktF0abVoTYZQtXRNojfV
jd29uEjfQtp0sSUDSfdAMSFqk/p+pCgdYjQb1PlJNE15hLqGJh+oLC1Il6/82jX/7DkXFfj/d31G
FSWVMMrgMicwyYCGI9q69kPHxFghr5RI7pvS+Cv/mtQfXgfBxZIVyzI8rkY1AOCTamsjVb1Lpw3O
jD9JFpHalXLD2iQpWT17i+lE8mqnT77iFbIvOjARtpMSa8Daeo65a8H+NFia2G2ij3h42JF6R+4+
szkscYJMndY3S5aYFt4xPRUVNYhnXN8/4kCyG8QIE7NwfYm5tQ6roIb4QZR/WF9xLCzILQk7eobk
c9xkfv3CPkiPXVLDPxBemVb3vvD6UWYSG8ECirtyOBU7WzmZg2aooTmxIroBw1X81m4uSpd/puhJ
YK3AFUb44wDI4RvGRaNjgjb9hXwtMt4B/dvHu3e62zkcpfDMEXKDFl+xpv6ExLavr3xXlV0Mps7E
XFsG+3mV5YOp92WzZj1VKq8GMuedjkueXNBLrr0YcZLC92zJ4JPdswsZWFhXvYi2b55GtYkC7M7t
ZX6Em0bG9KUYhpIPiaWjUnP46NNOR+sve44E62OUolFzigZPoOvDsf1AQ1Mkz3Dnwsopg8VFJf7z
YCqmIC8tMCM6EulLALuAnnp75m7olByLP+fK7Uy9vZJYvVWOBha7CVdRaPIosH/e4BUKwHmEHDYx
iBVJ4WIH/8VyUK9AUXKo9I8s/+dOU2xggpucrB0ZYdNGdDbzlFjgsd7cTDMs6TIHSdSUImcczoYv
GoL1Raxoyw3AfI43QfjTkwmI/S0GvRvyg/BK+vVr6XEgIhIQtUda0sBlEuCuL3KEXi8O6RH9NxBH
mJyrbyt59C5/vahoSWixXXnhXaOZxoFYDSGkkntycS/X+R71vcgUzosPcsMm1xJEIGzMff9eik7N
jbN2b1EnMvOgOqxpStU7MDYQbJH8/STCleGcuITmjwqO1UL6vNYBOs+fEH0KHhRZi/0THJwIgJOO
E7gHwfH/7d04uVoeCzePdzDG1Pn8Rw5kASQQK55/kxpJGw61B6wb9kDTHk/u5WK+OC4aUNnTppJ9
/3p3qmX2V+EclpgSaXc6lGpDWdVcPfRtkNG5y3zNUD6+255UPJBLeMcenbgsdMEdgKB7Hc3+I6WS
czqicROmaz9wf34ySOfr7AiOLPNu2XGhLFh5ZT0Ydm45xxlp4dJABMuUOB3m+kRuv4NQVZJFt2+x
7+1vJEXMuumVrS52hIDlz1w40lbjTjcedPts8vFvRLXf0hgKLyHi6w1kcI+4BGcndubA36DmfknL
MZ+S43pJHurOyOxuz3WWbrnu09YSLbHRBJ5BvEFxVGpnzLxaWBQWVGyrjP78ODxBxvrPc5rZOWXl
HKU0heUZbrptK+im/UZfmyd4PfcPgr5IPGn3x/kkEXAaTBx2jfm8hgex98kcOdSxgA8zFljgqQEd
y/DvjFmY5mMCmDvD6jTTJAcT19p91Ti1K1yTtGBtHgsWP/QdOEJJ9Lp7hTh3+pCP4oyV3Q8SfVWE
ACnfVzpEjLO2KdF/PfW/0Iiczfg9fKDZfeFo/EoadUuhnaokRL4aGC+gl8rPB4jIL201SCbUXKHK
u7SPUaIxFhnVClApKGX2pLvEbFISztix6IXJof+zovMUyLjTxPktrBvpwW87QzAF69jxE67FvoOy
0KoGYMZhwkN+89P/TJ6ar/0imPQldOYCJuttTq1N+t6dp2LtgL9y4nlPyynBrMThLxiEbdRqjELm
atbs/4YUWp2eXjdgkqiJzda2txaOyEzIwGSlWHLSh7xQWmcXBCazbNdWS1+nx7wBusIXGOC/itVt
uyWhdLZqUdzshpGlectWeDWMqE3DIgUjhyMArWjmcd8GvMuAJSzoGHnWzhGyPrGyTGzt5SC2KAQj
ccUhjP+r94eoGM2/t/i7dyPVXuJ0zHaWpvs0W4ZP0+TzOfDct/IOMX6bQem3x1n87sJZBdWC1tbi
QHZduc47q2JPVnezOJRmFThAud1Eg/7H4YyCgRLI4q7fcZe1NFPpqAs7l3SWXjxx8WPJkkv95DpR
icnZWbI9kHG40mi6B4y5jt7lPJwJVfBTxpjB2ZTkRPmQphKxApnzIolJuR5XtESdvf6ny7C9njSK
65Jr4vDzeGpaLWcuwBMAyQo56k1hpE2Qt76xfF5l4fbzUcs4HdpnJ8kKMfW/ZbTGbYacKVqMuMGq
6cNoEIE4koPDeGoho7ZWSSRFZWrymcI6fz40lOtxT5pvAli/6L+UOdFqvECA/zDzOlH8upgdxlSd
mt5yyBOmQzcQDrZ6kLpNB4lypB062mLJZtB+QNcbP6k2426AQd3d24krOEO7gYDXUUYxvO4dAMF0
xJLnHQhhUhkHf0Q2/1DyFn+qTwArNNicCI/qZteTv7bH0VVYT6hEa7wKkIYKhNeA09Wcf6g+2a8j
KA7Ad+Us5LPmubWq/Q0j9vapRc27KaJW41gph2E0niSF59UBatJ6gyVbN52n/MKa+CzEA7DvODJq
CVn+avP23kOB1bO8xwt4+MdH1MwnSMfUc1X2dU/eR4gUR0GzU5R6Asgl/miaAEWJo4QsR2BD8+z2
MmPNtBdplGoWaKahbn6AXKZjT9M4nHFaWPxogO3PJumC8ATGVxZU9E+54qqIGvGMYk+01M+VvljU
3jyGwSfrgC0iZYFH97ENfGYdMUU/n/ykO+FD/39r9UXA1xhLmnrrWFqDtfoRCECQX4rmus4wkDZb
x4ZglIvkmUAVM5RTBkXqRg1U5ojFqiEoz4giLJJhmPMKXs8ClBugPQ4EhbspcVvz/9nGCPkREo24
aof5eNkLyqG6aH4b6DUrF/o7er+WA8xWgANlfAkTRDqrKaBgRmzbHvzxpKW1a99hiwwXK5uSQ+25
LPZco8hmH+L/6o1yIgt/6lRQSeLklK9d7MDUMBu+mUIo+zek9Veb/JISkjL4UvXNQ6kKEk/Xvl6b
AQSCrKJEDeIvwQv44/GEq6Eny7jB6//MOq5h2daG6mE3bjgCC7DdGtonmG56wVeKneVKmbi2t8i7
no5GxmstrJtyaxu0ci8+hgbqE1ng+qp+koYiyFvjHPB89nZ3FdBzwQ6NOF8kpvMjwDGH5D0zAwKU
oSlxE9K0kgXRNT8Jvbw0KlYQe0Nsr5pN9WWmt3wnKA1PuEvr9Ca3xY3rGoQESyEFbaE9wM+9PUwr
kOjhYJ66t9++XzJ3DtfJyvtwboTrv2IXobSZ/I8JvT7JWzU/Eoc/Z2peJYtMLH4vB6LFPWL5igfE
pbjeHsT6ey10h3DizV99aa2ropK3PIFEhHX1EHBXvNxNNAOnkJmM9pefE5DvEvURAxfkF4aoPlp3
Blkhq3dFw2v0zh/izh0PAGzWzOZx70waX6MJrLQqCT0j/Jv0iE1zYdQOLxiV8o/Fnu812zOG9ix6
Ul7VUSXqnVTD0gLjX4NX7CdcAKYWjTnY70IWtcRbnKvJYKCk7Ts/HbiFrvwQNpTLUA9+tNTmzkhb
L31xFHPCopiOTmHTs49zuUfKFq0s0bLu2U9gDUSpO/Qq5TW4Tqv74gPRbltPvzaP4/Lrj4hgxqrP
OBoTQhiY/daV/7isqLbect9I2jmVd0UqZpd/xlHeq89anOf/gZHyCEaB7QwHvhff6TXrTCb9nzIQ
f+hskmPNms3lY5wUs8D/R+PdfQ4PQOXZSB2wysDHQOWMi08g8eCsL32g7Uc5wX18itUZH9AxMu4j
ysxjMTutdnI8er0gi6lmPOHkP5Dyr+7QsJz654LjHWdeZh8M99Z8PF10BUDGNX94yCHOFqM7fAjG
+2VlgPRBN6IBvbjq6uU7GijEsmkabJg5i9ebGlmZMGRsvFtvZK1KhHxAVzIk9Xv2ZM4WiiEH9A3b
ca9VOLUxZmoCgSngAzC5LiOqsEaxNZa3+sfRa61BK1drg2z4pPzhjmQFstzfsAwDYeIDQn2ZGFyS
TeTwim6dhkNhGmGNQ1mb9hihAqJMPMnjhPzgJq5H3hSZf/uhTsRxTIxg4Q/KAOFeIKjdHX+YnY4i
u8XYLX3Y9OUbJ+p39CYeHgjoILK0fizPW1wDv5Q+/NExw1QUd2W+6ShkS8wZeU1JV5onXCxJRVdB
kIXCbJhgXEC6xKojuTzRtBc3h3BQIzaVSRjY3vKacx6OJMN/OT0HC/f81spVUKKqt3WG7aoRvMgD
68vjaOYRI2Wn/pUSCRX0Xy4BFoJfjUrAUYhTASZ9lnWjY3rF40Y7K2BNpZogKsMK6NFqhnvqtGsN
eawNwuCB1o7FV9mYuagB+mXcoeQrsBvwpgQcE4PzVsYYgdZCDho7OFMBMCgRaiwMx8uFIFaIH/tr
HVkSr1FH6QmXN0Z/v6vLs7SdGIwlwjBZps1wEa6Qw68iBEpdmOCDq7zYA5eBRetECILIxu8jNllT
b+/SubwBP4QHBGI8oQ61l/02F2tRag0W+1ZETsJbuCQlJpOv1a0izuUiE1wt+FJsX2CXIcu87HSK
rTV1yZ2+Z/3UFVYcsD8U3QmQJjUjmFcuyMCaY1l7HVcpYauvC6DKsI4r/0jhWwSbMZyAH0VioK9/
3wfUexa9fGkrqgYIqGENTifKCE0z9wqiDi0dX2qmZd9MR3dRvffc9HmKItEFV7ycpPbmwEBUmSt9
zhCgIc1OGed7R2lIX2y7zhnYwZ7ixtQ5BRFqlIkYHMmOEcdpeyW4uVExiStNPXG1YzxTdB5vxLsx
rcsQf1uQMlb9u3hK0pyClmULFKLYB+zcPMVqIANuy6O0ZqMLff9eRBRWqJZSL4jXhhwdiq0NqbdP
beUM8EzEDG7biCmnyNhKPf/OxvCCIZc3p2SAy5+jG2vu+h+Pf1CII3FK18pSeg0HKzbe5r7o7WH0
AeGghwwuTLCoWNnPaLq33DyUBOjTfX2pbmLxCgyoVAMW/QWw0dv2cnmKO7vV6gtP5Rhv6cks1nXy
uXB++vJ7cZRlkopp/4Lhwv1rz5YsNEIXWSDml508/Po4RwljNdog1x2/4qks8UPbECgk4LSEUkbD
0op6GsMZP33aowXMliu85rkjNd69Qx7hpAFfvTYBxwy+d7E0y+B0mRDV4GWHw7x3DcdKWPHb4FHz
uACtfzcIw0ZjIZ9aE+hAd8WQFRGR3lvRlsr0FiQpAxH1s3XXt7JKf/ysLoCCxO7XQOjQwCc3ChH0
6ywAy8CbFwAA7kt6q12NLExBL5nimjb0hX4BumpwzB7v+FMWh+NgF3o8uQMQlPYVWfC4G/1z3Cd7
aiS1CBJSE7PWnq3wGRgcmaa7FcQ48gLe5k/12IdsfsDiL1RkGx9B4ZqevK7Iwh+lNDOAY70vLdBa
OfgpDn88UZ2eVbvwGEchV9kd2RY77VuOZ9HxBjYjm3NLSipvdPPo8WraQ90KNh/bYAGWk6/whu2K
1vnpaRTe6oETEAvXOtGxUvEvvspumGUNuI6i+/F9IY3Xh5hU0CD/f4g+ODi9pwoef2cCe6i+fv8I
yGFBEWOv3gOLNBFVf0cKZ2puY01Prb7alcy6ID8ABpjlujJc+YyabyCgC1Vu36iPdwJgRexgdlOl
ie3Mx7R1Y1JckWQrUH+9VZh33+tnkJ0sawtAhid6Vgqtfp1Kzyz31zFCsXMAybIlKHaMzKO2Wb00
6Co31oHjJNtJNhoFCgU8KVWLQz9p8hPsdOsyQ+zgRL3tl0Yl6BDMFVcaZDCiu8Eaagma8pydzCT1
3S/WxckGu+N/QaJ6i8Yj1X1n0764Wk9DQkgRZai1zHwTdkFzFC17U6QV5XpvSzuYrybQrDC17Dlt
DbM4NVEZ0vo48w7XR/fcShJhVr/Kll6zBYmNaxIxeEwOQT5hFtT1bf7bTwVkUPOI8oLzYmkNxapL
SzAfcJb0hHw5v3wmI95WcC0mnf9bmdEin0NM4gI9COig3wFrKbkna5BCPtuIvMiu4wjGl5idJhu0
iuGkDbNBxdBcOSRj+2RfOqFGn3ThJMzir6kXwmxnx2EeDLBJwZYe4ZUMH/vu1b6WjPdZ16OVIlD0
+qSbpTlHw8jVHV75XQ2KaSJbAmT3Q3ouUUUu+JjT8PXHvOYDfkbtU7cg42lrHlLmL7sp1YIuLqkr
qNXTf5k1sPSF6rtR5gkdTzCFuA0LWAnNM0+AsU8vjafwO7KDb0iclMpCYnLEW2IoIdlBytcsgQGo
3P12KVopUAGU4pC4liV17NwC13V+F2dvvvpnwas/5JN9zgo54UKJb6VHDp5NRAqIdwSSNzeYG5NS
j+L0yD1tgYN4V+4zPqdvVmx8MmEHo9GwM3XQFr70RPxhC8z/GEUf34S0afFJc2le44EZ3l+ouAOn
mOsII4fzdy6tQgMv248fGydXOXvS/HruEAl8ouaN9Uo7mVrC0+VqDtZTCZapdEmmMxpuho4VDeIw
D5T6Zm9ultUk9DKXjMDF/Cd13xsNc/VNrnH5EljaJkusHOg9Niv/YicbRemh+iKpePxFAo5TNYxw
pYPISQY7cUoWnaaDainH2/sUp3YveeWfdgeN2NbqgloxYMwAHwyYUkKm8rofSc1Pg134Cw8uPZOs
hSER0OT4jt44WrfwgT3yQyzjvd1oE7vyXEjJRHJGLyfZ+YGIxD1Df7mnKw3C06obNfsspMykFSl7
3gBDyLWs0fnK1sFXoUbpHFx0NT+bbMwJC6iL4BxRmlsJ8tvkrDomx0p7wv+66apTuEsI01kqKPJp
en7sD67vG+uhSf44BSaVqp2Ep9Epzb72JvKDo4+5EUObbVXiRGokJCpftQgCfbikR6+/8qc8HqoF
tIyU/O5/tZQAzdo0OmcwalDeihYnbymCdQZy/mIEbTqxpaNxdWupmG8cjjv3xqe17S6ch/WhXmHB
p9PEuq3H2OlZyLjZ1CM9ow0naWvdp9YRUdPgY/AUTAgKoQxmWq5NCENO8EIPhnQJ1wLo3X02lWyO
axGEPsDDE7PCBDAuu+Ld+yheJXa6CPOa+965H3r2SGjD3vf/bjcqR84lPW2Bm1isn/oxjTXD7lU+
Tp1MEiiNsUVVeGmeITiX+HVUgSKqSZUq+uHh7e9l2S+9nh2ZGInqM9G7W+bkv7mJt5xdcTMedjMC
iesbvcjkRto+Sh7IfidKbQus+kgWYxsd6n984ajALuyPALRA79puA74nXmLSofDyNJuQUCXZadvq
g7HN+0y+XItDyoeNEseYJnOQTO24ncnvak6uqlLEkWg/ZzOJRkjzGBB8wyTYI8SZNx6OBxwRTCBL
wnS2k28B54W+TPkK3tVrDPQc7APK3pIylHlN0qoAn3a+a8U/n7dqsnRt6ODRlvPP0x8Pt8xVeFu4
5bVbM3V6vyjyWueKTFF1UKrNURT36s8toGaZNC641Elt3FD71jmRAoPndQZfJosYle2d/y6G6EnE
LVKinmyLRyX5eG0K25dsDc3YVWsfD02tnVK0P/y6cqNSMHOQQfWoos8julHSnbI/V7lgnyN++wWc
Nq23x0rAQIjvLUiRGl43BuaDst+mXRR1eV4DSeLuWS0+0o1WtVD+yRKcWpYvOeg6ODFs11J8vvEi
GrfAOxsiJjJKh6XwsvdNq9McbQ1ngVL6ezYogecjS4DqbNPZfx2bUsFqCerhMBojCIZYnFfkxtZD
XfgwUpEMI3Z1wgyeRRR/SjiJUKBfOfdVsifdlzkfe72RaRYD7bOSQUvdieEhol40X6LhayLKZqV7
VeHe4Nke/UhDlTHOy58IEus+GyD76kQYNzgE/rmy6pX5dFQzPz+UyTfrI2fbn3Y4P2NMof2W2LWz
d6zT8ZVga7ohn16qxvtv8Wf2pPUy+6pvlM4fF2fjQpcvAXSHYXZ/ty4ZRgaekVQbTlKaR6pLbZr2
Y3AFX2hC+GgWioODBxcE6IB8IJpDAjkFBvRDJiH0ClatKm4/iGeIIl+AM2h1neR66u5AquxGGYp9
gDSCwodiyEzsdJyh3d4Dwb7DAhAxfqHbu2enYLoL891bxge8kUKdSX3x5E+aEjLMs6btQk/jNUag
kioI5Rpd468dL8INXYWzkQZN8iuYIATi+ZxnzBxGk0zPDSsQe+QSCFTNArZyZI7rfC88SZM+A4Ms
ipUbr8XuDowfBsziIdG+r90cpR49pz9MtjxaYbAituyhmaB03Kvvy8mGjDNuF55PsO4yt7wVEgm+
NlRfKSZEeKDXsrFe6KUV0Jpg5R/Rz8Vz9NatDmmAsP3Tg2qPsQYR2+i7uRq/aC7ivyJmhTzqHI+F
9wy4djnLnmfrSywRunWIIKFms1dW/zgITRCWaAsIGvHClNkaZGjSBMZqGLbnacrdkkIU07Pz++Kx
fZ2Ffzx9lmReqJJkiiAo3V315w4T1rdFkqCYNMwnonL/FYJ/a03yFjQeRiDn80RYt+erGxuUs5bo
LeJQm92oEc5uvRgaDWWTgZbHEI+lIVU9fhwSGavmFE7iFRYETYlfreZGezGPKuQULv6S9DzFSv7e
9gRC9D9SwD3oreUq46Uh4d2RlSnXcunSZaM5lhCEMXcHkvztJ3adcDqDxT0z7ag/PrHfc9l6DCpw
PG0OSdFn6AeR7pBvRRftw0Hv58NsAr0vagmoATbYBsMc5/vv+1t3FUi9cAICyVNFv+7ZDJkxaqGc
oJmDWRthpEKXqrGG9PprHz7+qGqrS9zApliHIw1K1kZtbH6xFhwZNeg8MIZjg/77D3ecmmGMfjVW
9Q7vqEVIocgRSOqsJPKCgzNEDMf5ojuwPOmlLv7ys7y51+1sorIfX/vatH9ry1a/dZIzvLAOXVi1
pdHV2G/ZVlOx4/BENYTnN/nicf5D7kEdbKgyEBlJizxl2j0tRcxOV5gWNc41awycM2tJMp4aa4SX
mtb71u46nSoVrBmQMa9pCN2WQWQjfBekHjDspYUa+eLo8rsGibq+mT47RCckrvV5NNxNKJbbxt0C
wCePeYZB0AgnUnNpYJaL6dhW4A03EGrofTU3BPk2EoKgRz7i4K3BVqj6uxkyLCJQYQ339Cie6y/T
NGJyjeTMQLFz89X0vk2BvzN3XL6uiWBeG8tSplxAB/3iE6T9s75PyuapilFmk8xF4RzhueGcy6sd
kcs7m9EmO4ryCHnzx8Li3HA3AfPRWFkug8WeDVwOM628CO38OgMprvyRABGQBICwN1dTiAIEkpqv
z3uWh15tVpMJZfe9NDkZeKlOL4AKAkSJ/W6QWj6Y86HpLguOOdxFurWgY0s81urnlS9upygZbrZx
nyxN53gF51e8xjJPRKoJE4fqcvaydC6ficMLMPjCUcaJUQhUhP1ErwkdcDHNMiv7w/kenz9g6sCz
a5VWGvkhBUWEhztdzwlNbeduGc4oscV+XyeDip+vq2u0Ye718xA4rSMOLifsVpGt0FvjIB+Ue617
58Yd67U+07QMtKaSI89w1NvWC+0jONz20LPgDQzwMBdN/UGfZjTUEmksnk0ygQNx47KmmGp8eocM
qZpu+XvjZF0ayOATGxofO+1WdoiMo7nV6dFV1w/0VXwr4QelkNRZo3jq2VLj+PtjipPs/uASDdOa
6DTbR5825W7hQtzeXI7EhUOuKpEvMzGZg/+vg7P6gwVihKBuw/Xl45Ock/MfSRiKiPaSwhX1P9Fp
3pRHdqhymOfcpcUKTn61nz8nmcGLlPTcxx3mGEHkUju/OIhUxAusqz/tlNYubrYCF61AH7kzU7r9
TD6tq0cNmuAI74gVaxdAhF0mNtUoaA7dv5uQ1go8MA5H0CVakexZM6CipGHxL/mV7N9QrlLZ+E1o
weD5tsz/3xkwfr8wdv0S5GLHJbURtcy/anYemazgTy5Bck+dS6SenpJLnkuRs8u66UMdITHFpSWb
R8goadN/4aiEGUxJz5dyilJH0pteCERSs73DM2nTFapFb+RI55d12VdEOjWhYa346AoCbfS+Wfff
71mXdObo+U72ZZWkUQpewkH+vu4HK5ruM5cgj6KqOfvaTW0rGcQ3pqFCOQB7KUaftazWsxpnSsai
QvPP50ocjgoy84fCnN2Nw92kSnwis6dCAiDgh8NpPZpQZ76ywim+GxWfJqHTHzeV1P/Js2/BiAHy
4HQnP60Cqe98tDO5rcpDrDsjXCt7H7QVz1z+VQbc7tvJ1Qw4iW7RYfjvwUNgRfwAgdHCwCDZfA+x
2WGdioXi5gZEyW8EBpNoLeew3T/za6HG6Zg4RTzUhv6Z38fZqWO67ekZIUB+fNLyTqd4IKRpBsCe
H4/60Mn8+/1Aduh65oJe7s8Ro8KK+gJ+ANH3jAE7qvPBYZhR6zjnMIVHjdlOt1SWJ/ay3geX9LBT
xownt0xjmpivHrB+C2E7RjJjzL5wfuzSjJhl93n6Nv+YRVcybGuuROUrK3cj5u1Nu/9dZAyzvyg+
XZghJyn5RCLOIgEONb2bi0K2Xy0BQeVj1erh+5QKaa//mg0XypTfGO478jj0XUEBGKqqvf1Hvp76
dFsSwlp8VfwOsdzUbhfzZnm18CRoAq7gVE9Q4Ch9ArE5xg22TPlJemlfHP8ewZUegRqdogA/+qW6
xGFDCoOTlALhXTu/XrBpxwoC8crwF+BkrXtmEiRG1OY8L/W/YDNUKajrpiO/A0bjqGgqfe8mLxmE
mbenZgzhTLcVPCri1SUEutOlaLDPdXLIx3dW8p41trajnO3dqlkU9z7rFcfkLfBO2UoIlfRveplu
xLzozW/MzIerYE8whzaBa1UFPrh5KudsMTm6+nrL2JEYQBWU6xUyiQ56VA4gQkeIHz82ma02jkAY
ZOUXu4oT+o8i3sqONNYxz7qhBtxw3TOFxzQoJqjWiiupLCdCU3p5g8MAYT9FYqke/Rg7aCBukJwQ
bETp5e05sP1SN9ufbo5RS7P/dn+XgCTQ/iKziyVVAL20mW0UFWFenEhi2l3wiesGL/b4QJRcbwv1
b13RADF5qNHUrd5Kj0FLPbsjgqCU+4B/8FveyoY3z2Iz6C92O/5qgyOcqf/9i45u5gwokJQn5saf
/FQNJW9fSMAAhqu9A9rI0Wz0ejdf5WM0CkiNOzyDkWHim8bDIxyEo5BHtBcnso8m6f/A3V/As9Lg
kbSEp5+nePg97kpr9OusgbcuG4ZGeqPUAsgK0HpI+cx6kfM/F/E9M28nQssxOLOj5SGdXcIzFMw1
ezdV9YboPzV2khPlSyaTTfRiHfE4PpTzF45QV/z9ohzZuZEoUd8YK1OyrCaUcu/mmq/Bxj2V2kbq
xav69CvvxBnglNyt7Ju99inb8QK89NHf6xgLU5b4z+Ed9QkXuktrEL1u8eOZImsUWGwW7YUJ5Irm
THDjM6ySpXIMTZiGIbRf1dbLL0RTspMeNrrxl+1eMD4o8Zh0RNRl6PxFWxGoA0qLM8B6aIAH1IAZ
JZzpmw+MgeBQXV+HeyQJxeptV32CTOptblJJxPlCW0zfh6kc2J82aaPkHfXft7BTBBU1jrUuLF5H
i8dAJOv6bD55hr6+K/9zj7PTE4t0iEg15CumWR8i0VGTw2ve2NTXh9BSeR0NAimhGvOTEbYTgsNu
s0QJcyHc5wb18IU+6PJJSeSWG1xNQY9qkr2vhffCRW08VbWp3VfxeDQCX2Gp7ecL+ttDkndjulqk
QJ3otsxZXUo/gUzAiCLoLo/A9KjiTldGomPiqu2/tRbwbxsx2SXP5BK034iF0r9Bz1xtDlny9Ls7
mPKV4zhEj/QH/U7N3DuTVFrf+zBhSe6y5rpncC4XL/w4FtPTgbaEo+WFI8Ekw8vGdZsN6fOigUON
W6eoUUNBN8/CpbBbRDNxd3tWBLmTjPNjuZZOun1z1oRLgoAGdWZp1oC6wQKn/zDCzpKwhlrqL73T
2nL1maEgeI9ni4xVLT5EyNGCSKn0O+9/sLQDbtzmEA/XD+hL0wQD6SgNaVS4IFaEweVY07UhrScU
ElWRvKbIrofUozydmy12gLcXfWz3Z03enRfRsB72LKKA2+Ev63OHfg4sn1i8Cxb2AVz7YxPSoR4r
glNArYllc7QYw9Ba/aH9wGM+/QKOVRsDtuoFM07Ad2eEeJEwj6EiUPO4ai802YCVgALxMrxDv9SO
uhSqrfHWmNSMMhYPlbbhF4osFcz0BcpWv8l43Rmih0v0K3MZiDoSKKxwyqAd0LtP44v3w2GEpscP
eZTfd/1Zpw9irZJTALqhd4PLbYkO+dsxQHqdorS8XviqN3k4n2iTKrw1BbrI+lk3NNj9Qrkx95Li
1b2pBbhy/ketdUkLNZFgpvV1NwCn/MCpwTv7t2bw+el2b9mnbjRZUXK4uLgzsJ/85Ppk0JHWH42v
NDuIlZKWvtS9zCIDlhC0rUzeYa4XKdgbB2KuqHcy1KE23oJkjiNk6BLCQj490iPf97ZOTXfYhwLs
2G1w9mIfGGK3D29OEVrpUkGvOc8VUmXrFAMG6MZF8KDNzSUfHq6uJTdXASGAb2GorZFApC4exmQL
6YTo48d+V28bSZ1Ol7/5ZPr7mcx98/PeJzb5VZM9l+qL1DyBdzOtpGbhZEDsqjeskPV2aCjksDDI
+KbgILp3faIyw2m9MXTNOnTIgPw5ogibp36TCzVePAarN7xw5bYTlNMzPz21eNoye6bWE4GNy/qy
sJSMAZKGe/k9RtgPcKQ7qsk0ncQ856GcvL/igu3P2HUPgppQGQWAgmWB/2J2QMweDtWQ192KeKEu
omtiSR2LS62VMDFUGzLFZz+w+WTMaEm0Gbs7Opocw5Dz0r7inoL9hNvK9zSx/8HoMojYKGrksako
49TP79GnGOkMVOOX0iXhdISiPK/hAqfFMH602CEmoExVtD9LseHsZwHsk71L/NpK9w7JWX/0zgnt
D8LEwoHAKIdD+pLamyWd692mHY1mwZOQI+v38ghcXQpYb+JIO2GlgwogWSc6esfcvdkAoMRlScqj
oPcXizRz8BMr+a8xWNoxZ3vJKspeLbs8OPPvrObSkqj1nhvQ667eImNXvl0wNKjZn6pT28gzTXlO
3ARap7BIvQCfMQps4sbo1vmKu/RWj/QtHzX13Ht4t1xsE9XKysZzu2ZUR81p0oH2In52EAHbzfgJ
LNjCAxs7MGe+mpJ2B0ULMOKanlwz/wmAnLbPLxluEn6e5bpSKQTWpTLHdvSQnECya5EgHVieAePt
QMkikrjNRAdds8TS1s99OVkxxxSJMyx6kBZMXHZYBiItQjk0LWAYOqE9BE5kfrn7696FqfCgiGkb
GynaQc2nRXvB16I9h17ZMCi6QmqFGF8bvmYapE7fGyYUAtQCTZ/J6EtbT/8wH+T45zkth+Nh925+
UGP/vTh15EOoBOE6RK0h4YAzOFzlJ5y7sg/ehpkL+pRi1maBs5UnsvCemI2ntx92oVmc2PEG/QGk
Ys5R/kXOG3pVHck/23ztyapA5vxU526BlO7rh3jHvNGIdkSnn/jelBLdTXo7ka0XakHv4X6wPdA8
RkvN7edHUw8GUTk0yP76OGfkByiv9+Hz2OMkjLhpD1zbKEGY1kgBZ50h+DHSdyaPGXedwENvFtBP
7EwBnV+dCt37r0krLk61A6OChn11GQBkBd0cvhhv5/xCNiPsrK9Uk0EobLKWLAgloJuWTGezuDxQ
TJxxTdc1DhSOw3qzUD6CvWo9pPLsJSTJEFeQHWrim9fNZHkIdT25amlwt2pae04vFxHwM3FrqjFm
+aSJDt+djqvoPJOfELV4JzKgf6/24XTT+D9c6IKGG6iOqBfoDtzeTajIlB14EbqPAJP++SrJa57Y
hw6qskAe1+odZHLsmRihcT4jg/qkQMvqEAWdrLDT8DSsU9gLE0QI5Ruw+8SQHO4t7LKci6Ne0PZz
c+8t4i/4POJxo9gtvhdr1xphFxegfaZ9tS+owBvf/yfdpvZ+fxgvDPI4rLf3us/XRWWw8Gr6B/a3
1OdqXikPfbWoEZClsY0+L5gCz7wV9fdVPKobtdQhesuHvhOSOupZeaMrrMXZeavFofMOVjK2Yj86
Oa10YbpvWLYD4wEc+GiOGU3xNCFqjo8tRrWaeYgJuysVfi41AeRg4WQ6kRiur4fFFCBUZ0h7uO3f
DtNOvo4OFUy4O0X7hbqlDdf4t63mZ7cZ2Vs3u9bmWTIgKsTzNTNeyeUjhdtM3e0udLW3h/rPEUl5
nQl6bioMPlgxZOTHQqCYOe9bRDrWZDoaOINJA8SsZ/+7RXIRh7jnO1iLgskDRPSXGcLiLi6dqzWn
paHMefH1aKkVKmZIW/BcTFpen60KlDUJ5HhGIQp/EzN/luNaKts/kOEgX5v7wp65yxLi6NLmlzmh
gSF2iHxQ8uYCtoV03Pw0E2VR5IDTjXcMQUALQ0ykUKGJZnHCZGxG2nfnGjxyZUg/CscrzpIC5wxT
eG8xwA5GhL5/RJnH+ZXQHIMyjDlhL/Ow/4eNVYzGSEiMX707+20CkMT8qb+7Is4uEGRg/t/vYWlB
2FYvOwYYEQ9KWa83ectxnpuFC344y9z1IB6cPfA8SyCRW1obYoox5/nmb3MA391t9bYN3twdDUkL
z29xt/hKsJ8uGkKQBMpe1QbwexschFR4EL+lucR53RT4/WSu/8fdYYs8LJ8IWKUDp2SWgMt/i+tW
ytzP4trfrreG8fBpwxLhzIGf6Dn425kiKeUirU/oIBUoJAegiTQ4l/UmnvRtHZA6MTu/ePz3wx7R
0kq3Q2xPSHnYj2lBmyzuT9R/rY3K3vUELKzWxQPO3+FbUeArJJtqVBCd85WLUL/4DdBflXEBpC4X
KBeTKKD1l0tLE7yR+JFgkB2BXlN0ebYbCOsHa0GRAVOZhBoXWyq6rALjruWJzMQbnLiuUL3pbl34
D9o7KnFUQKDjqToodKZ0k6e9y1GPGt8vlOYNXy98yxg9B2o3MD5Rm6jbAdZfueHOqmvoHUyCInnn
+FQy1GD3Lx80vf/0RXm2Al+RMKAhhbkYFelDXg9kGHJE3vT59tEj3frnlA7RYkJF3gP4zXLgYG+I
B35O2dnveDaB1NFdZ+lHZWl5XjWeeFaLdJChvodUPtrCPMDHuu8Kb2VpjwyGJPnBVZ3jCBv3otX9
vbRhCAuVcqOH9kLXR3pEcg3jWjuIUWtlnfl2eDtaG741DNOtQbkEj2Jv2SV/hw5JSy5QsdVb5CWt
LOTtBL8IEUrKTgx1bURaNLKvj1M5V0KtTZadm/XVM+4K+fK9nMTx20a1koSADzI1Nh7OhUJSqFp+
4JHzZsjrhyCxrnEu54pwp1yXuIZ4xPPQWUdALUGjMoqebvRNb0FlGwUJTjNfOoxEzbg2o2koGUC9
BDZFfHCo5Xfgm14IQW+gXZydA4cEZ6zGceSZ2/KotndaMx6micarYdPqzJtYrBWrWoSNIKajJn5m
ws43Gstrbnd7/HbzIBuYuekPR56B6Wm97QROOkhpixe4gpJdBym/e47vYgjFpfeL+uXHM9TaxHUQ
bUcrenAg7j8Fq3ZCuDRVF/As8pRJjNxKxH0ql5w3qhHufohjeUerK+rX1hOvGTSQA/8ND2q6gBf+
aACGYeZBPd11gGftJ/5tgOlaArp6GFduEGlJFzW+upjsgn5ac+ugnJwnqX8pzUBsoL+4Bhm61WWx
wYeeytZz8WXP4N0SttJXQ9HHHdYf2jKJs5On3OdrASfvBAGEk5uDEIWwMGl8JRpbsLE1R7ZL1PLI
oNBSCjNfMqIh38KCzQbl9k6fks2J68+mtmTTYwllTIGQhBeGh+n6bsTIi/iEk7FaDQlV5Nb5E6U5
gFQHYI5B61Oj11Jb3S/nwGHa4l9cbvt9TwWwINfZZkvlpKcN4VgnkID0yV6HqK8doSjncYmq2oa1
qaVg1xKPJFyFWYiwfeeX7z/ul77UA2GRlRDshg7C7ypwFqaex/gg0ybx5MNpw/KPy5yQ3B0In5il
DR10syZ8Q3SFeHVxe2qndf3x9phGh5yZkt9FN44R1zgQhOtM5eJSLrYvov4/DQKXo/cCHE2lryA7
5AkrZBc2e+BcMcQF8UzMHhgiK+AZZJKwu/zH74nFA56dKTaKFu3RL7BRCMHgJBh1s2ZOx1A2LVIL
yvonE38oJ+AbANmoyXOnUumhDevuZGqqmoB+9ic4V5YDsyexed9vFkPR2BcSVT7N9942bpyzFqvm
FLoWxo5m3ZNxPZ1rA5UMFiCHJQTNg0mT0kPoFbGzZAoNxqdWhOASpSI79JBBKt5RBHtC/j3RuDS0
hV6dehXq4OumvAt3uypvBS3f8L7MPtuFu2f7kJcseYGAQljYgyJkrN/mjyE5Zip0xaI8I9PshKOm
N+gdbhfaiQ/l1ivNXWQUd8sTkAB9l06sAi7+BKKZTa5W1aohgyYCb7CtIrWBs51FeqZneNp+PMrD
xMIyeztFdtJEy27FwlyZdeRP6mk0K8BzXh7p1tePwseqU7ivKrtLwVS3q9nMKk1AbwZCja+AQ44p
WJFsp8u9/efNqZghDuDAThg3ufg0iXkzbfD5upzFYw8bZfkIzg7YG+E12VtmsLC7zfrpsV2Xe+8C
/kHv0IbGhGCacxC55/8B+s7RP1MvTO4KDOkumDdgb5YkSn+LofkhVN2SYgZATcIYHHJHxgv9TJaz
G50knfe1mxkRbfQh5wTe4UU54UFwN9r9pufWvVqv4MgLArEbeZA4b83Rro88ydrq/+oNGGixQXaR
GyxexiCxSvbQH3wMG9EUrO2ef+5RaoGq0ltwIwhhQfDDt4X1YX36vUht75qwGz6w60o9ZAdaEfLn
Ceaz10F7lGS/qXKRjTY5PzTE6sUsBcpcIiresNXq9zT11z8cALjGr1+29dqNg0SZv3OVFGvDhI7y
/eNJiTuKYu91OuGMPa0PjnnRi2nDb0H4dhvk+QA9YIBOjviC+7+R/Fyk+Ji+5Cy8X8sVZNWEI1Vu
NfnJW/Rs2WHMe1HAZViiTvsoPu77ljN4odwszTFoXlVVrNa6GIZqsiti6okGGpip49ox2NfcWT7p
WSiqnwrsKz0CDS0HqiJSnoezhTL/qdfsTMEEU4dBOKL7hody1pkP+VcJuF1eKj1ftWnz2WqAXclm
R3vE7aoErvaQaBs+c4ARmZL9VMgTTT0jX+wRVIPqJdDR8QePombU3AygkKHaZpPvvh9AHdrkkIVI
W/KdBrCIQLvFfL53Mv5ay581wdynZuCyGbDbYC+FnhSMPy3SOc/wWU/q1+zowsTFEYPYbrvY3/z5
4RNdZvqYTXzRdpoDxC0VqD3fgR2zxuQu+opFwmLuCHRe24G5jC2zhhXDBbxtt3mi9vhSIX6YWkfc
cYEGfRmae5fTqPJMjP56lngnCHQAilZJc0BT7U0jxvvmsq1AORT3i1dArIQ7uHcH8T5vH4e7Ygji
P3TbjROjI76ByWWJQG8BrB+ovHrg/0EUuMtFdnfcMe6Vb1cnXjCpsKeyr9n12l6C4IkxwxsHvyNK
6LxRvXxHlTsDFRMseG8YQ7LdSpJ0RrZ2i0sQbTThiFfnVNEE5J4fwi6oXnFonue8QiLf5KPVCL8k
OxY+sgnh7sbjv/U6oxstLZnJkH6Mc/BQ2JpOOiyN2o2fjoPvdKj6//NF2BKOkaHLlhFkIoJm1IvL
M27tCDXrm/r7Pv9qj2Beqnxya179a23HjzmMP1t1yEovLIQYO+176bONKl6u4yFKaDBFW26s6tDE
snL10bRT9QbUmnpi9DmQbhJWXHe3+HbmvfI1rL8dCF2XyeaasOxGSYw0570fwP9yOAsmsf1wbBuC
g43wlDMp1aCb9ZA6bRTgOuYj+/mwZ+8htuYvJkfze31+zHSqGxJ/YN6bVXIHjFh7sGUbOXwpXQaj
rpsbykm1mJ1p3VZFYZqm7BrbZLxvtr4ESJGgH6TDshc1BJLDRUlkMyhAjuXpEgaG3rErq1PpLRNv
Tmhs+cxF4cL5VFY9dBarfZW+u41j61KHO9bKnNYycUF3aeLyIvsrq3By5EHX065qs3G5mz4gdtaw
gNO7NIl0zHjbW5kU9LRC8TnNGoU1JktPIVUW1rw3ZNLzgJzuPjh71bm2cMNc6UhctBtWcgFpp91k
+y2SoeUaj78JamK/dp2orihKZIgPdhHFrHDquuN3FM20rla2mR5ek5SvoBdPakI/udkSCoeU+DQj
xD+pa1kUlYvY8geKn6nQqvVcUhpTvXytfS8qExLRFbHPLYeae8yRomikx2Qta4x6poJNBMEFJU+G
0qfrejZMLqS3OXkHII+Lk5yp1YCgeszcBX3ncAaHYDNJ4sciJpngWRjqCnmpz9K/uCJeN+ZkNep6
JjXoasW6hNd+NWmsPWrrJwIXbv/7VPkpzkjPnmGYNUsNAlbL6PCiUWOjCRchfr3Fi150aI14qmzU
IQhWEMbjOt8Q+y8GRlH3m6KjweHMxJ28/pEXwJnRrPUT0mHs2ACjH1CEVpisDa9X1iqamCYcI1wn
xjHM8hwmGycIFpO24zTEPvRbF1c9XVe4yNVZteCAV+KGlRH+feKVl7nwEYZhjmMkftGp5G8ihE4k
qSCOv6eMraxD4mm18WUMoXDRjF1is6RpvxrIcHphlsqncqZZpElKa7b58H3JBypf0FXd7kipuE75
nzfIHaKv0GwSxsB64poost5zmlxUfz+n8mZurIPltCjjSJ9x4MIh98Cee6ZWLgLhgjwlJgUjYdwn
rC7fKZhhKKHEsjeIU07QaYHkeQgTTWdEqRw3mcmm+pTALsSgjLr/NukqPzTpCjI1WgX0+y0UZP5G
Y/Kf74SrLlqytCjYE7JFRVm17WLFtnDxsSsXl0z/XcePoZNGbnsk8BYembpjMSuWwqjnnh+w4iSP
tOJoIivKNA0mUufWIqXvLaoeYg3zWp3TKiytpLF1kStjJmiIJuBnNcVgypoDUKXPwcx9v68SwQbc
R9obmhtsdRVy2kPS2nPxRyTDfvd/WGSELQRGO2ywuK2EDzKqWDld/lobZ/4SMas9FRiyyytjdMre
ITdxoTifmwmUrLkB8OX5jL7rz6knoOAXGM2O4p/JbfczsKe4pw6KG4ixkAdIa/EB0IiVFBXEodU8
zzGl6obVYEKWsqn4Mu1NgMITFeM2tMps5+i/5rA6/GH02y8MLYfncPX48tq/uwC3M41QmSOv0UTQ
QFtdJyfyKRmSZEs//KiDf2AiwnmVvneR//zjg0wRTFqViLxUNAun2WvE2MMoFcqAYgNMcssVabav
SNLkQlHJaLSYOqrOPwxCEHE75hEOUrgtUkIIur8UwBfNujgLuVJQCcAtKhwioiYqmT1AFvffR1tr
IdBJ+lutLAzZmvyKTxBawOkh230u/p313u5kQHRXj9xbB42DIMf4ccp2yHpH1ZTvIpbraOLW9bMR
lnser8PFqlETd4fhJ8KvdhkMfjGTOdPjHWyO8A0nwpplSL+tiAJXUjn5WXtruN9lBlVbfTXBWqip
mxtAj48h0VOQDqTJJD5FkuOQE3JjpC+7eMJqJ/CuJFpo1f4+m1QZDti+11AIiZegf4G13wtz5sHg
1LE2w+fTaXaEfa/rDw81rHVROUxnZmqElur3fm0JtF9wT+ZLok5uaY7PYsG7Lx+B/tt+MnybuKI8
xUgtBfy2RZGPt99e0l1kFsCckU5wWBjc03Oxv8DdAfnC0d+RXnPuS4e+Z2y05kKoE3DxjYhJJ021
AO4fvoLQYTsP/70s2QHFy0XcgEdf2PbzaiHm6a9mbKObm1754tYGSyFg/G771A4aZJbP4uOp7aSy
3VtElLYbWKXU32DtIedJq3kv/dK+LCOX8UsR5SdBpCZ0nD4aRsdzdAZDpMwfdMfnK/IYOVjmGyXX
f9cbUJKAenpYQObufmCNS6jXGN8R8BYAjt+0SrspUHL051Si8aW40h+x0H1PMDxVeMACZOxuoqiJ
Gm6VNHpN4LCFg5GiFj9udLGI1N/jQtKWXUqJUKJU2iVNtnN7kzqNV6XQHvc2kT/T2vWpw8E7xJr/
VVAEiZNdD782IvFJPKeXRiazhMDyrpF4QJNdfcPaDYJj7MZOcorBhoZzl+4l3NIhynsbqxGnEbUr
Lexpj4xdvblTccs2APUWWRexDzhSl6PwdOwVxJti6hdKcRda1lB9LzYFo9fkbWUv2bZyylqS8XZU
3MkX75hktIEBRSGawHrsx9lCMkmgkSNEX+6ioxcanvwHy5aROvH1PiXWLwmFvxVLoHUijrQ0gYOX
joNtLEssw6sa1c4MMQoaF4Qn4/KX44abGFa1hfpghtSPgKgVLPMLjmX2rOej3KbjC+t2oLsmDc/2
ris/dJSTlEIicewiq4JTgyUSq9rsZeUrDvL7oGax37LEEw5CEkWEOsod2A1kw0BmAUITY3LeBRbj
/txDhhi/UeiL8LWUmoBp5H2lAdTFxx4cyx5ckSyhzAOFZ+om5kBREbv+B6HN/JVe1T9pAarcy2it
HbXJ9v1siJOj3xSVy/ra42fDLMaBiehP8i5R9ZrMs5cIBFS7Bor8ycIxODumhSbAN2WQFOpDwyte
QRr2OGKMzD3zOvXYVI4lg676V77QKgQYfiiakwQ7W4XctQ/GXT20phdS3WPzL8Gy5rleJOpzxWHt
0mAzcmSUiD8ga42lVcVj/1o16RMmajdM6XaXjXI5Nhh4/kMVAS19bREyfX93PugRRCA1s790IJSe
j8fpBsCMnRzKgQjeOPi9cKqQQa42RM2cyApsqT1kYTorTqB8SbwqsSp/2UsxzPDRkMkHNS1cpWwq
SvzONXCqHPjMYo0OxWzdF9zAUdoL9c96hNzwfxvxwSmgi/SA9QvfkJcc8g3FRIrdhlVc9pZ1cJMk
XYryGGfO82sTdR+q6TLrZ9rG4Ly6JfkNYRugUz9Iy01K+rps/qjKxCfmOE5dyki+O4mlovvZD6uD
jfXQW1stXU/euF+bpLQicQfAJOLAloWPdKIL7kDMF+h1/MQyKvQeH9EztuI3sZhVGPAThbjpR63H
bfgAW9U4/apwDF5GmfD9gkMRjlphW0IreBwbIgKv3Cb5n59xgp12VBz8CtXlMnaJD8kew+MeNxP9
KZmpszgBnBKlXCnN9KAICMBG8blM1smaY0zpmK/DtGSR7OXeAWPK90Rw8JEz53T1mxo17B1fgeDy
dwbp1e+pDt9DVRDhRXqwQ3sbtRWN0qUANpPH8dir24hQ5eEuuEAUDIb+pWnbF1pv3iuOxTYfLLsM
3UpxzGhauzIQYe1kaRXFI8t9EExVVP+bggU8r/pTzhW4fvkkjVPsNxUSvEYc8hYku9OcMUxmEbzz
efBPLArU+2PHQ6tds+coB3X6YKz4o9BCuSOL4Auy/6LxjSunVA9135gh8T7tSwyP2hTYF1eydGWY
qw+slkIgQ/7oJRxABqWOAdZisnZMCXT4YDzbjgr4RCkvlrj0O+jDq3AstIAMsUj9K7ar3w/4HzYU
3uh7oYzZioT/Pn/6rXwelqWL9w4Pte6EtOXf7R5QhJAXBnQ41gd6Ud1M7O2XU9k+cI9zQcoE9+z3
80FDvdLbn8qc3cSu8XzBG9Qn0kGMIg/zqCLBUNSC3pNAptjmgMvg6JC4U3PKqCNM7cHjT2e0eLre
71rD1rswkM6Irmo8R9uyypvM3B5XcUehpLNBzwk3GBA4z/Hdm7VoZ1EQ+nO5gcFwCUjtVMkQERER
mFJE/Ya8QO9k+4QyXF28vA5D/+9Lg9fl2z/Ic8VRcGcAOSC9UYvc3fNm2T3Cr8XkwnD45+HLNvSH
lV6W0OCxbICcUXMMVTb55wb/jbMctgjz0vl/H8PphVCdAg39g35bQnPay/9T9l9J5RLKKL9DP0y0
cFY8o3BUf8WclaR+ElzodF+w7ypXC0X8M2TiJSKQUIuMOKZ+btoKMPx98okd1VQzvyPBvXWniTu+
DYXsFpe/KvW8FWfIVbvRbwMaNHVrkl+bA1SruPwh7S/RR/rb3crq9kbVe9cpxLlpE7LCiXBFYeKM
IIVGoErigMxzdf4nZwWdGpvefdDGVw8IFqGREE3Jd0nJg5zgzk9io4c0ZFN2HJrOLJtXmmdA+SF8
k7MzU4n9+j+ECwb9TweGjmyheALPen64nt5deIA443fD852xOrRFnT0zBEqznJecEJ3YQf5y3f9O
MJ5shak+DDNF7YeTFt5cyispXnI+uNPoI9tNvqKsstc71ciCfmPTh6SiJbM2Hn2adxFqLzyfmL8B
sQVHcIT+SVp04R48wFTReXrpjGjDtI2HHGapf/3uOhGMzwd8lYrmR2XH8cdy7ycBxKEnDNRfT5DO
XfKQu7Jc3PYu6tRzuMDfy7RH9iUxNFQUEIqGzUxeTe6OEtzfU2WCt5HN4GTB2l/qbP00VsPewLYJ
ZVIlHR0xvWiRQqX3qfKMTZHruleMmQ0zzVc7ccQ80Tl4FhQiEGJhQ5uivi5L3pW1G587Sa5TIAoI
FnLVcGgMWJWe2hLOxjF8k9PSkB3xb3zSig3sCrp4d2lI64o4SMFV7OucJZe0gOAnCsh+6DUJE0xl
zJ1HyVX057156EJ2SZqkys2qDNWLFyPRS+eyktOsin88loeZvED4H0K8GvV+GMW/4OBcP0YCdGuS
t9DgzgqjWrgZSF3MX2G5TSL2eyD0f0FCFUAEqek/bA37NIoLzGI8n5WNjBp6DOn1+GXA91VgeZ4C
JRljvrzbAYPqNW6HEasexl4w/gOh+m3JkLjHTZTuMuVVN0LxK7/sgXjjDT+EbzMdD7fVkCQmhnmj
vJraVEKGpDKB48ndXsyhDscb9asBFf41Hf9h1Y9fddqVk1mjX+npkjN9+AAR3j0WD7SDu2YmXx3E
ioKCFBpRlhjtg0Sg9CLW72HxS2G/8RqmtRFJfpeD6gxpgMJ/D/kahXt4w0B+FKuv+UECjdyJelzk
wxA2Ps7qyPRkyt1GM4ZFu4aAclV2ky/rvssAN8N6hFdO5GKE5prOTsftPsspS4frRCP2SN2fYntM
Aj1PGkFmrcYcbp44bKY8CoLXBs8FztXMdPc64wZ9rePi2UZZDwq0H8yTtLML9Vgz2lHor28tyHXd
9hPsX2pKyGT56e2ez3ipo+x5dFVJXzJVR54RMG2DhNERhjNmEj1XogGt6VYPp7Rxlk0T144g4cew
dvtBMFVxtfDYKSWp5OD7WPv0+EbWhw4QjdLjWtWaoXH1EZbU1JF0AJfgeSpTVpmkrfRoWUHQg33v
gIjR9JctTfNbtPaxvj+ouXP+vnOwB0OcNWrAUR0TJnh3GJyCbbWf7LDLT2Vd0JxA0QA5SPtbauY2
wHzpl+L1s/4dYhF1xFfPxZfs4IlYfHPCgfs5GFRiyxQe/rb1CfiDNMEV/UEzOSlvd1vMBxV95jXS
caDGNpRL4C2AqevPmPkH+X2LF3ujEp2JuWzLqT+y0aAUW1DoBnP+2d8Dt11NaBYO/zP65rF+csOt
CTExz9TJ2NNmL/eveopx2nd+4atARP+xP158Ur722/7cRzreHMa1D5W31MwAoS+j4T8nrFj1mA1p
vbTWI+VPgclFCrD3MVXqGRARsLQ4JKzvks8PVWM09tBgMJAxt+BxJO8kLEiyvDicYl+CHpWyP1e6
PnCxqrzcerqCZ4pABuu7EtdfL0Z1YWkno2/Whha0qoEPCk+97B3S1nUZZLITwMnq9kfiz1TWlGyb
Es5dXPcCCPBwYIb1GowPn8okq83aUWiUbl6CAqF7cbhLJtuIdhAvbSqDpNc2qsWp7TFOrU/UaEAu
Nk14IPP8TsjLX8ss2+85X20Y0ibSDVAvNIyxFYnbpUly6foqtq+RXMNCnzbFRlvIemm5hLvJHJQ7
lVkIt8smFbW+U6BtKxlhuZvGnMGWOXNn8W/QPkU2dk/J6yFEiFz0dpNOpfkkqspeIPlku4A7Yz+S
qTWtKNjkoKNJlCm47VjxaItK7FRvjfz7C/hBCbyZDco+1vEJz0yIDnUtTbgCY5DeArVGW2vAh9MA
Ui51XQnpY8wVqmxa3TfkESvYsBG9A4FrX5LIAHdvFCrebtSoOBxVjKEImQmU2TaYZo6vCpbgiWVX
V0ZDMTV00sDcGYpSBiFhxiaW9GW9i/yBW+sOM4jtNdDx0vOFdY0PoXC2lXWmMx8r1sey2CfnjS4w
yDxaypiYdxeNYfv9kTODmbZ1ukd83DDgKLqPehkenXbhMpMkeXZQ109RQn6kXLWpWFvH28Pujhfj
4YbHnB/Pw8BSDTH3ib6UM9BZDof9rtBmBT0oe9SJUhhXUn0/4phdKzBvy5M9x8Xl+ABHQt4ez/rD
KLvaMCv4niDq391WUQwqTsEMAKPZlHEbKeI45gRfObriVR3bV2K4TnUKKcWlWrFkOCM1n4/TQnOD
oHXBbSOYOzyl2Sl942Veu4e8Kmq+4ahdgcYkDX5Q8UFHblVNYkhJibQHmjTD9o7PAcM1rhDzeOLp
LzbQLs6F8El1DDqemRWrMYxROhQ0z0S+PDWjcQUgOLiFRdOFg9gpDyQHNpFzfZZW3tw0A/RKKZ1B
TathnqrV8jOFO7UqVOEdcFYe+f5w5q0AvxGTbp7IzEyoJUrg36VJWVugF/HXyAF4G44ucemeFeM4
11VRNwDVZyiZWGEO61zL5WXJYEPKyB7A6bq9kmZqY4b0GfykUz6TYc7ta50gByY7mqfZSSe4v+Ye
z6kKZBrbSzZpEBhLAaKUV8vYdL1SCCMX6vqr6agABD6T0cdQvOndco69+mw66t0E6YnWtgdQVULJ
wYeLprAdH3le0f855UBvzWjbJpXu8b0vIz5b7auKVcvMBDtVfmdbOaGznj4f/ywOhQ3rpPnGYfTL
TBCG2OqNL3LQRyV0wddiLoyv26D4SbyDh+W6P5ZSO7rDUPg1I9lR42zI+rKhJZ6joIA8JsDpIj+m
GozyIK0Ry3uxO7E08VHzZ3e272jNyxrzmggOB8yrHYN3cl7Pt05Hc4mdDX3askfVYbnUm5uZR/XE
3YU/2ChflKoe70vvG89ODwlySCDuVp/Gt9YrImupfxAlele+25sOXF9a/03FZhupSOPxUmSZjRqB
WiHXwt8R3hANOuJMeCJP8LxnyLEjSQRch+abRhpllflmLtNZrJTghfeHcXiPPbAqWN2Gk5+0ciXk
O05RIt8Qh5zhKAQClDbA/bV7WG7R+7A8TrbrZ61p8wn5Mg0hTaYnWUcijPnuFOqpZjbbp9P5iskD
PAmBfFNgzTaQEvZQdPcXJjAJxw62d094w9mmEhbjWugS9zFL8m5t52OCHZyD7NSsPyYu6mzizPUr
amqiQLsXeyMhXirxBNvFIDllEJh0Kx85ulZlmhsbQu7FtO4qOWSNo0C5OE8AOTlgojz3Cx8tY6CB
ERvySHRT3kPm+y22GocmyWtUK9BxAySMTEDvaq9gy+VJ6lMk8qaO7rtt0PHN4FFYs8zP2mUj5Hs8
JH/78ftx/KGFh8f3UNr8KQ0DjLDuBS4jDpjyVW9tUC609bqjIUTeCSDyLkMImClvsam9enmPtYI5
CW/28NwNMY4rlnLpBwUNyifJT4ssaF++F0V2RALVDk3lkWGrQLSoat/5ZbMrqpARefTVK7w3ffIf
ucpY9eJP0WGJfvtNcIcfKqMnVL3iUiRAIMycnhoPp6QZsZq3GLfRQiTYLe4MByPspTSd/eZR0mb2
9yU8ijF+cE/2fml/3Ibk627GfbRv/GBR/yZQ7xfiq2IOKGhi9JmD4xZoB+1cXzucwezKpoT1f+8V
MwPsPH0SNGhLzNm2appajaReI9iQ7Tb47lxTI16MYqjZoQdoBfVgFEt1lnBfuFpUAMrmqMvZ9DFY
UZQFC4y5VFBVSEPiVZ9hjSxhKT2Fci/ORETzQf6yN5cjumZYVuFghyI/ou/aarRYwHR1VgxWK1u4
Jot/jVGpvJFbYOTNiER33qZ14VPcMcXHEDpxkCFwFAkrczUm07FfXChe0HoCAZJEEA5zESvtr1Dm
E1895vN+tbJKIuhk5yLp9UNhoZb6gNsPRJEUSZESvRJHmJeMFPLieFYItnPlWmpmt4Z9Wd8PH/vW
hM0OMbO6XF9JTksB6mGM9LQ9hmFJgsw8k3rGVduDxuNwTQfSmx+zl/8TJbdEyegg3vkbCy/U+YDg
IutgaLyol7qUkZxgwzv0uofK3zHoLANbPTvZzW7Dr5GE5goT6vo1HLR7mOUXlAUxXjOs7MCeVZWB
BAV7RbkmwpoOa9/+sIGJGjVp5+7jeC/R5O0AIrZzqc9SUIHPrKJdUO22+BDDjSyhUNvuPfvbhies
bjRlvz2ha2tI0hviNYd4DVGRAszBi5c2epRpG8tkDwvtEQ33yR0yrU7TojWPV/84HyCutgQqcAFO
cBnR/3iGnikd2G5CHfnUG48y+vxA9aCbHBH0WtUxw1lylfJoYEtm1+Vc/qhXEPfbwUab8kkiN6W3
nrM/R206w64i4L3IK2g4oZGzVp+b0w/Iy5dNrYRompJIAj8Ql64KtfPh16BGLZ3aYVobPQGzxWUG
Ix5kPfqQ2lHex8cv8IAK1dJyh5iiv4B3KECJwTlc7i7MlPhFp9KcFT1m1OntH22cD2n3GP8bIgTA
QH5C4BA+MG6SNFp02CX/AytRiVvGAmfh8Oy41+T+jvf7+OdMG+uPKmrJXrVJIf4jiwfa03b7M/sV
XXeM/GnTVx8iISy+Abxy3yEZzsk4PuAqoW6VwDv90xvu7OwmFkb8Zac+xGPvc0IqeEiPWw7mpHGk
+74nSVG41QX7a2uiElpjnkYiswsR5rf/8Ln9pZr/UnyIeNKDTMPSsjxaYo2Hyai4ViLbrQyXGDA3
ueaF9OHkPt2zKx9KKQByYisG64ByrIV5emG/xTW8Q5QzbJWjJHzjxpVHXEE+lkZOteLdBzZ6rDa2
4jzp1SdychGBNY3Q1Kkb7/+W2tGoGYwX5/5eTNbQtusTRyCaZLUKF9bzNS3o7ZyzTkPtkb9xkptI
dmeIm8QizOfpNr9zpC2h1djbtEl3QF+2MrNDwW39P0kUsVP/oqOwGsndg00pXx5mHSN/xxizekC3
XJtaJM4jkDJ+HCjkjUE6zgKADBWjy2Ffn3gvWWp67g6zJMCkbRN7Gr+hk1BizZYJN1Mzzo3Ea98d
phs0NCBJkxu45KC0oqCFvty0K89bJmNvMid2qgJ6FWba4aaryBnK+nqOYJdkWgtFZv96GztMNnIj
SGLyoA5BSsEIAVmrKTO1PWbKZKMsRXs09YMuVxLOE19SQnoKIe92jIVT5D0CCFOFNVY+0yJQ2Vcm
t86nKbPJSxw9l/rDLhoQqO/Z5dnmrcU08kgBjU2LmsdT2V41I/byTMUh1ow8zjVAyTQuTI1B1VCQ
SpYArYXG9BEI36MhJXjjApMgG5nJnujly5+WIC9OBFAr8rD3iYyJc8+Vk0hgGa3XXqBPn3bO1zFy
iR2k8JFrs/GGQRXdziej70d92No5hPdcNgD4QxZwBVbADVzQBQb9AX0W3STog31yiqTkh2QA8pp1
T3+isLD0+sJhclhniHKTfPW+WmCbbnEpYDMLCEWvw6YwEAH/yNJkDjNZTLC/jwNrOIg1qZVHNn/z
aoWrcd4xPh0t/TQrpXmsfa0MWVQvE8T9p5vkG6TSJXncIqtWZ0JUIQhKzLyn1u/3gpUobv2uZtaj
4P11gWG50QnzDszVaVW331uW5iyfIpPBzxRjiTqrWuDFB3J1eiUKtzFjnaBVn8YS5JowwU+WWPDc
fbwwRkjmALefTaDzmW60dBpYmrE5/SAXXFurklOQBPCZM5DDIPYFfEaETKsIghpU+naxYij0SXDr
oel11yfh6MevZ5aFwEvZaXKQz/3zgejfNIqdybjz5+azTe7z8pti/LR6yhSSRsGVN+dbZljmfhAJ
jdWJxy1jxaXNJuOfxDv7u/EIFkU9MTHRdOfqkPHE7O+xHFozka/SKCNOiVDMY3HO4Ezk9NEWLOtK
RUqJCeTf06Cwt8JsCKmgAOtYpfybrf0w4o64MFvr3h37lfV6XTImINy/9tR0w2BC1Rr2B7avBha5
iz+2bg4ouhcgfFE+TjGiygAy+nFo9gmlk5v3TTuaPqM5pP1d1cAD8XOKw3L+saShs3w7DRNtPkIT
xZvKIIoNm9UWWdL8syaJ3h4ZWHBw6fIKQfWyuy0DIsnN45XZtC444nbi+JivL7usr+jPJSV3z2ay
sIrPIJ71ckSCBZRr36gAzE7GvcMQXoumRBM8k1WlJMCMQg/HzyomgxunS7HOMhG9v+ORFdOUgVRa
PlvLZiSARN+XcYEUDYJXh7ZnRinHSUYgH0scELfZugBR2U0xzA5UZiWKi7Gr2x9zHOMyrjOY8o8V
v8PmosFlkxR/hwxL3EVhNcJorysA71jQOWq57/gGzzfb4GnnFC9qWUpt8fZHQAJ6kqhJl7oz+4PR
Z47793RosAbgQ8gAVlglv/nDFhrvXRk301nbhtTGWDRy6J+7Jkd1PmFF86i+kF3UDJNDScC6OTia
jlUHirbwe3WwiNwrIiG35+ZHHslkju1RPp7wMiQC29rRYVcOpQW343iu4cOBj8vC6JHbRt4mqF6P
GvswiZ5AFjQkQ5mZhvxHtTwB9Xh5fUkmNud4F3Len/iMQLAriT2cDg3sTYD8qCILcWxaYQmq4TmA
/7TnIyXmzWrgR4wqZnXZybtsmIC6AdCf/ONqZP/vOKbe32SYm9mKdTXuDLtFsz6R5wvvGhtQrUHI
nPWm2m1Z/BDuC+95Y5QxSUCF6dkJleEEp5WjgBoToJKNIqsqyp1hA4twroeslDruVIQL9KmvUY2m
a5geXKuhDigVlD9vvjeNfUmm+Iup7Jiv+6Ew4HuCEVtNd1QiA4b9Athou772g+pwpesxkk9GCS1O
DYT8XAIojdi47ETF03lGOYYZ7dF4bUcN4NsMQdwSUKlWD1DU5vXdbdG2JYPL9Ei9lKHcFy0DTzM9
u13IZknGj/SOuFQkE8e6ZtIJKvNIS5AyA2qRvupxZsJmIlwI2ffx7VEe9ad01UWn+IT5SXJWa8by
n01haupf2Yf5i+hIhmUazY478+ksSUxLcXfOVU3qalGqtxYjEdZMkIZ0YBb1zMA24pKb15bXyG1d
bBExCfvASvYZVRY8ZhXw31tTb6G6k77pzt5L2vfg5DkKD/PGgYR494Mfu/L1AYV07Hd4UAvEbhBF
LkpquJZB80aBAC3Zl6jukK8lOh19pGgJ6ebihDQpTKTdkkE8esd/chzzk8Yl5IJ6QwibxnPv2ZQk
IaZmAHiUwK1TbJNEyIbMTuKiBS+ffXPxpxyPWinrMWHdS17P5lQ9w5WYRJ4AJVYNzZUYnPdpJnJV
xiLOf8L/8az9PUd0cZU8srmJenAMgMxGq8TmOwX1IehvXgUi1JGaD+iHkLu57JOBaWVAw4EFaXZr
TcrmhOwkBazxKk0DgFhtusgM7cfSsnlFOlp6eFwWPJ7c2lVkAgDcL/HowBAhf9QT/kqlw+wkefP0
yCy5NXPg+X0zRd8XQQMbQ+pW3trjA3XB7P8E7KTsK+36UYqlDhDucnNfc7Ifr/7lpK8/KxHMo5fy
iQFGitmNS8cxIiYOdlk3tsqu1GfSIfZtgqG9eqFMFRzMsX/os0yE/cHiRPVZE5qjRSNJC9fIYrFr
piRIiS7fAX14vFWu7tBuD2MC5TbjWVvHa+CpvZGX7reTVQbHWu2HhxSCk0xcddxUesQHEDcig3VI
ecNCQoKjbLb6EDUpCwG21ZJB7qK2HVhMcEuVrRqVp2atJ0i0NSbUF8oCiAHv2mV6QNTkFWtmFfXd
/GcpFkJ5/m9djlntEtLAigSSctkkVRvEIFSX97z/A89mmkLrKQppZO534zh/4VYTovgIPx/qg85d
vUwSF1hc9MaA8cSiSShlWLwLVVgDQ8OS9ZBCYSw4Z4Hb6Mz86FD4tYQBoKK/5YB53kNP0UFB5RMP
TUqXZ4iRAohJzgqyCcodVGbt7LC1u0OFFy8dMngAms8kFcbZYzfbu9zwltjuQ98Htmr/vFtXdf6Y
bNhgcTnOOQudAjXdLnOEoCfmq6lIkEi5eo/WkADTtN1hOusd7DacDEsLurboLXFbUBFsCuxk30Df
vNV4/H01iEjjHXbAJyHfuNEfYnvxLcX+Jkjhf6OB0IQUPAdPWxrW7tdvB2s36v9RDXI2DqoiMLc6
LKVJU+ceZEN8dTJjjh01wLsKhuNr8BsvDOYvqYbnm6kaxezOM1X7g65kI8/E3QB+TncHoHDY9mfy
odFTycmB5to8qPfrcBwmEsBjX+k2LKYoCaFDRpzPtwtUuIQCN9zX+4CowObGkBuG75As8f3SD2rv
vp4BXuv9pUDlFlofMaeeAE5bMZNDa47F/asA3YXKzMplyXU5raAT1OlnuCdtt4I2Yt4aLAo/xNjU
ZsdHyPbkWkVa9XYGWl9IohVsgOcFM67t0iREAwqWLDA6ad4dQgpNV6DZpclQmO71WrEy4p+cTzvQ
2a+KyUO95CcSmj3Ry0EZVCXjMa2E5oY7DDm1FqbDxP6Ug6hJpC65djwd7qTijANmoCPuSMdMpQJT
DkF9kpwerCnA6XbYBZZzQIkb7CW7EG9IGiO/CtBaaP7wCdt2lvUG3nkuLXDkCoK9q97XAa+Q7Pr2
HLKUe8x6hRiCIhQ8SyUS9eYvgc26KIc8qnVYAYNDS+99AhD9D8vIlEBA90EQT6cmVAWy7Zzvz/rm
iL0iPsiCFP+NVdY0C7gC4/hy2g5OGLqoxdhtDfNdxT+OtQyMYU5A5WWgT+t34Hi/1qxArrFwlJYM
1TYp9udfcDMdyttigDa2zbcayMA6y5hTuPi874P4kBvg2buVSJ722ndXGeEMqZC9DPShMfHTLbfF
txZtg7BlDPuby2KTbRMj6VtC0yDf8L9zD6LjxCEjBnDCig4pvUj7yjMpXjzYqzN8wQykozT9ys93
HHV30JbWMeP88jh2czxG3pL+t68H/98WQHlBIyuPIuqhw1JvGnPoJv4btLI1/l27DPZPB+e/G68S
6Xq39Xva4ySewJHZC3SWUoXy4C2Z6CnA+fP+Q+yfZMP78ugTt1QX3KG6BhrVZze0onrTO2bkJs4r
SfeECPqX9ihWZYDiXEgmu5WoLja6BDa2QzJbwP1CgbS2QiPhoFccVYJ8BKTYTTikgZE4vBNES3hq
WxQxdHCs0I3nFVh+Iyzk9GVOSRzI1SCg3G58SL/3q5kujmmv8u69KvnphUCCt4ImUuW3arm7vLQl
US5aE8peso6XYCMHpFfP+Q4S4ipghT9H/aws+VnujC/FQ3yDx/GQxhdAmdbzYB17ohqQo5JEFTiM
EmEVViVhUY3ENTWXwkoytmdu7avktwYC9qVNOddJmNzL80CGQPjxbATQd6IefNDL6WrlpTdegcS3
oDKPDU3zHLEobdBULoBRiqtjmmVsZRJ6Z7VHomInw75CkF+WyX6i6RNOSp6u71ebYe+FsrNyV417
o224kEdcBCl7f+BsX0Yv3Fp8bMtb1kviFPVsQJk/qDxGlUibSrvydPWY8YDuUnlwGd9jYa1wnhcC
xw0+pBGyfN8ZEnVXxPoNFXFQV8N/nuJ1cA7ZuuHIWV1wIJvTyiG8m5/IzYzv3zKi8MRmrunZL8Te
4ZuMN3RBe0SyXlV+RK3p54S7JyrNDRvjlCTX4GHwBD6X3T3QTCv80sj2Ac1mNjbv4mn6MiDHMJHQ
X8+Q7akunZ4qsF4NQKOVNm7dh6T3+8dBJ78EEvQhWWwjF6LVLAIowzbIB6EmoSne2JePl2Lwan4W
sD+SVNyV2ADuVe7WiWqpIyrwBlwUy9Qi9Gg1PcoK5fktPuo02F5kFgj6mznFPLx1luFYjvOWXR+z
X9upEdMtTklAm9atDkQyU3zc3DdFkhkH20Vn1q0MlKxlfAJ3Zys2WS4QF+OHYjnMv7Qp8NriaGlv
DubN+n+LXpr6YMciJoHguRTuOrCPtwf0gaGHpQjaUVo9MUAEFEyX4LXkhcZvmLJoxJHflbX296Js
SgQhMmH2hR9Aq2Y9kHdWQTWcPioT0KXTA4Cxn/9biBDIXFZuCznoBinA/+MEWsasoQO3s777yf4Y
VVlDRHGB1LQzvCW3VCM3E/igmEYVJ+EjAu7vBSTYofnlzMX2iBjEdWCMgTykPkDUl8N7XxZQxF1b
9nRmeE4hxABg96IMxDQok5juZStlJywdd5vxj+0c7rz1pblKcwH925lkpWVCsgTRBdSB3iuJAHwz
PBTuCeoa/WI7ZHGB/IFItujDE+qCkhEAEKIY9S+qgPtjSq6mo5Fk0E8DjOhSbVixtPforOnCu16U
bJbxdozft8I2iMgXDf9FUl5jAINv2y23ekFvU6s+aIt1MojRJcmgZs/Fd79Cfs07vE0Qt+1YDHeQ
amTxtKiAnzB10ySVvO8sNDIn6JqYYaE57goolMVoloiQ2JHtktHeDCY2w7HWeFy2GtlDKKBal6y+
88v2gRdEwAeb1MlnI2bKs4aNaLDi+91QbRVPIIrgDlL3CkXGkX60qi2KULKZrpJ36zaw8WPvDgDl
hGUzWppES+yIQiNmySzARpKb07ljINuzeX5BMwPQMdwqb500m66ooih1Kh6fBv61hbsbGzEg6F+i
kDJNUsuDoJEhAhlIrTgaS+vQgIvxyWqH3ghB+x/mT41mfbeWfTXrMIbpfiJLh5eaUfsqaJEuvNb9
diAJ+ICpK5y1P44rjEOn3eZOKScZwzOuqXtxzC/O2HPpoqiy2UIOKvxQ+J+OQlQ/HVo0P9D/SU55
t0ytlabXFebkCy/RXCB5a4WMA8Adhj+igSdOzTo8I0t3HgnJsXKOJfygw0aYyQxUPh77SGLVS4R4
ZCZNkRFNSRv0sh8TO4havgElJj8d6GYvzJkTCosHmaULZxvl4MRoROJhHPOqJzwbttQQbcs1xGCT
1/VX6B4/yYEIchEEIFAnLwFbVtwHqmlMJOBUoRfI/teWB0BK6/L90QpzbyuxdDWsGNp59TYzry43
Dy/f3BTpgHD0+P8gU6o1SiR22E6P58jv303pTO/fgMMtgv4AVnBWmCXhldTMAkCEUqCDr4AzmUvq
hJ1o0C20FFANJrsSFV1gIi4TYdanMaN6vDWHfUVwL7YOHvGo3f30kf07KRzpNRGMVRWDec71EbC6
IwekLl6B6DQ6kjZPQGLsIA3Du053toH002NCMN/vo2WWNxscR7A46g9/x+h6UvN2PU8q5mg4j/Gq
Vh/O5qvdHkdDX509Ra0LsOn5KKni4s/q2CXqU5lmkEX+9+ADpcfTX6Yu1wnk5MJV/D8xpYg9+GaZ
YmOYWkx3JxaeAxVofNjgI+EUdeWUIVk8G+Y+jt0Q/1jZr35H8CQBQK+BXIV/3HdXCS7HuQj0T6X9
W7uJcxHSo9L+Qb/nKAxDmnYASGbrCVCIjQgv9tpBpMXGUj3SyWMn1QykvF0GL/GfDhqgxDq9SdlB
SbA40vpoFbmuV9TW+Se6mrCGPEmRrJFIT8I1K4GqwyEtQQ6qizwPMqNbJuGpwRKe96pr0+yjVkiH
J5XrzGmNZoPQ8FcjLJuf87xEkOXnwMEpJX9R54fiiE5/odQV3aSwdo5CoApScHSd01IUMcvzhS0O
LePfFqhxO/Um/IywU2sZXtz2kVJIjXRZevov5EFpWM1lMWueP0h0IFsM4FpOH3jitZZZD+Q8sRDr
KovTX9p+CufAzQGUZPRxCRy5cFYLJzYTwtLLn7xON68AwFwlnfJwigFa5VbzlGdFGgOoAZytysKN
CdMKAmUrwHlYCTVM1YdK3SoMa6Wzgc2niXh0LLgSzgco4MX8LQoZIeRlHoUkMTdbBb3MzbLChGvI
lyF5Zlu0rH6C+SdDjPqQXPvC80CXfl1DLdUXEIoIVc0wbFuxNWOJlQ/3Qm7s2TaduvadMBneRUfJ
iYWyu2rWs5VbE4qlKPf8nZf3nRuXlRhGXMXWZLA4yf9xROCuWT/S0wvQyDwDRWR3W7LtktpuLJEL
jZaTY2W/bM0gjSj8DGJkBYIChJS82xAjsvjR1wV/zbvXfeAWcWwpMleBZMt7uxllQ8pqKgNgYNGm
oLDksRUINTTJEZT9oHQAOP3sLFhNCRK82TaiA9MX00axFCdDLCXHugSFBUDgiaZG/Cf2icOKt99J
LSsyyF6xhe7AdaPYZz4C9oXqzi5cfViqTRgtDRUiRWxiJAX3eK1dZLvApg9ICrC7C7veE+3qV5vI
9Wxc3RLEuwikk3Is2qR8tYGTt11ilKhFcYYU5x6ZDmACNy+ulcRShpilTkmhA7D+rJnpj5OfYm38
YWN5T+Ol0IPU2rxVha1mXEqUYw2DG5Tg0SfHIzzRzFukFMtR2f4ALfiuawDlqn9uEv4lK1YzLk01
6aq3C/fjNLQ+weghX135yx/e7mErzxgASjXctpDT4hPmOP2biSrBGHjdJOmgvvTulZVm4gE4d0In
KVTHaB3u82HPgSMKPhWDHSlJhBofDU6on+h1rm3nZP3YIhHVZugftwXtpc02Gm1AfmPDGc8TJgu3
1lVWvnG1ZLWIDy/Ylrl2ErxLaERdKVhYGQb+665YsgtwRdpIhhqBgKq10WVwhhJh/ka/1cSbow0/
wIs+rj4AK13KUpR80EVPh7kmmgBV9uYi4TH6TbXb9h8XyAtB3jzKpVh6C27O+BG9Jf2WV5maOb/W
QrMOAXsCXpU5ZW4lN8JD9CyAACUR41uI82tVFX4Y/Gn8X+UL3dPNWWjLgTR3xZT5Oa1mjmmUGKaD
tmTRgqlyOafpg0AiYydbaySSflmQAPCIZNXp0PMOMkWbNi2z1GJRR1rZyS5ZevcyNcjWpONi7iYT
IQ31Xpg59TEMu/Nn5cyy2fUHpQW6nEPFQgqkz7p7xgXjdIzwMYJ4r8nCpUW1A7WAOdI1eJlhnlUK
unPwXzTCKhgLk+vCDLsgg+xQF4F987v0rReBZrEb/xu2KKX2AFFg0y8EX0dhomwh83e1gd30VISh
dMuYyW+we5kG1/QPRUaaJP6iYiJhJ4WkiKn7U7q61o8FpiNOf8R9WT0nLTjQu4RQlCTZwpLxESF/
+gICbfKG3P8/ggvjpacfF19JRVFQ5+gMcdmJkRnD37zMvpf4AfanAxmQyL5zgE7+ex4qnTbDStLC
u6EElpSwFDM52qNcLzcTnbfVL4MA40JwIpzcQw+mrj59cw0EIIrZaOLds7eDDdirgcHbN7d30fsP
oMBCtY0v+yCv8imS/mnBjqRfpnGiuprgvY3+ggcyez4KxYQGnKv3lnzwfTs5kZOtUtpbbp8ML/DD
Rnh7bnTVRLJYDpb/2YhGAH5QjoRD/fHxFyqdYyyLJxlIwtNtcnXQMg2Rzh7pWx3I4nY8T6nFLXhb
xr51xr/OE2t3xcKKVbytK1SxCE/uuYuGxG/3fb6vuEptLI85ByGuADN4S9JlUTjE70/DklzGk9S4
Dzzwk0TGuhvGstnSih+CufBSam8QEl4s5B3e+wID3zSTHnxdmsYlrrOiooC0jZHq/3P47xMkr3Vp
mZyHaLEq7FfE2DsoZOMdR0Dfqi6hSEa5Y1QJUsA3BEMwq+vKINZbUgGLHao5vCf+lHLpo/HIJr6j
/IyZ9aINFUJDhqEF2SOygaDxULenwD0A0RhnxzVbwJSVEh7+LIDqIJJXbqUJnf7AgmxGh2kUhnb1
5Ga8nzTbjf+wxusvm2gB6gaIfJqfcSTJF5j1XTU9C1SPePSZkxMYOYzj1gpoQCgb56kl9WqNV6Mi
8t9WgwmzTOmqt7hzFO0rfOZLb1/WbpEZ+RlCkqCORLPMPohMtmRdiEdkidVK/BOwILXVtdL5mOvM
sjUEidHAm2q+zlZx9f/9f+iKxNhRSxmVYE6uZt1AP7dsIsrki/nWMXWe9KcSAavpfborXxoPXhMy
0NTtOrvEcTuUcnRyOIsduwGYlcFJa4UEqo6p8/O6RZK0XR3EUTc5G95rIySbEuNVTG9VupkyAJqU
M20tlnnQraHjow9nE9q9IGNB0Ot0NSRNvRlLybNfC+438V0qBGooTryW6iWFiFKqsIO3octeWO5d
Tt3HYGOpZ5SloCvKvdevecbIBWb4VT3eRCzFIAaL3sYuZAjEmggSHu1c70JP9hlc6hwdRu6QXzad
4B8ynvBnljHToNe/ozOoYW3ohnXoNbOVGvZsXKYU36xvewQ5U5XY0EcWbWa0JEp6+aAcH76Dk2Av
56v9yeE2j8PikRK+3uvGD3maL2ZsvLkB4zdG0IAA4YI0fpXgeWwshpkG2yEnh4aaciQ2CaYiyEQM
i/Bm1iQxS5bunsceglFWLSSJJAWRSEVjyMkPb+6sj/wOHspBXyDSD1nvrHjdDgZswsmCRGDfVwe4
u1pgF5WS5RJnHNPB+7nAzludgLoYWf0eJ285VkttolzOeBKbN4sQWjrs1Y3bkC6Qh4ZXNbzu8irJ
Vkpr8iiMywAYoukUstIYICKsybzuk4/SjB8+jS9yjW3pcG5GOPjCUhmIGlA7Pto/4eMOHyMkgKjv
9jCXtm9nSyqU6bx4bbNMJXVhZ1XwKg2/ZHvkt3wvNBZ2tiEyBGE+vNXFlNWaFhK5TEF+3P2ldYLZ
oLvRbf7fSPb52A50NQtJY0IzwndGHy9Z1LUxPaeOcy0Qt3yl8BxcNocoaJ6GV4ZRlnSqjforUPjx
5Ft4dOgwuT9P+/MunthQCI3NYBtHgN+hBIpqSEzzXOxkjzgXwbaky/RDDySOf7r7UukLdzA9vOcB
EqW7DpLYSt55l6y5P8ebKiq1zSlyHAHLX7ujXH9cyMpbcaRsaIGAapBrdlxsEdqPBey9T0ILE5Dx
K4aa6dRmnvqkBy2yc4kxbfNjV4JkRy8OT23hiJqfjzwcOvkmCUlVtriprFXNiVU7WyIWfvCAW084
jSQLAOzrL6BTq/ECVTxNpcaUxDJMzrGzTObWxLtqoVw/0T0nHoYhhxcOWUF7gz439oP8Zyrld2zb
EWqjxdAN6VmMtLe/ekZDmL6d0DRcMn751avwtJIGi6RwkMFLUmUYqoOOAd6nixdxS3iUqi1M71BY
7mQRkYx7gqXJZBJVQ7NceY/SWUFWKaSQCIithjLGOywTWVWwp2drxwiZ/L5w4ug8zRiAmFj3HdzL
jDjS2ezgKfcv/FFDk1z2VQCF3driKepUgMQ9EpJmpYNPM+OcmJUI8aO3R4zvSrcKEU0SOVYY8mjx
6EH9HcklWcGT2fQwHet5R8GwdAbLBXlLu/+ixr3Gw7jOekKAs3wTglsLCuoOeNH3m1Nl3qtpJvbK
H+s2ZU9TCY+aDtn7GfETek1d2Z8tPtECBDNqfvrq/lvZvPyHD347x9JQhu69OdCCfNgp35gdOR9R
emrzE6rH2jpB5AhY0ionybupP1bVJhnD/p8z2UnKNGUJGFr8iXdk34X0iaJvINZZCrCQ6Czv5VnF
g7tfye1edo/miJrIXEzG4KvQPDQbKj+rWlK1t/wXmIgxj/pHCbqZnNgUstiJRe/911JNb2lGEey3
ydtmBu7SVpLWHZC/xqvaWF7a1CSDJrHso5cBhq3NiEKnRl4Jx56Qncv+OcMlJjklojD61F8pL3bG
SzAm++TV4PnXaeB6iIclFR+xEKiYODy2WM6N65IFaYeKmwQCdor9cmy6Y/YRMVw4SwK+uoyR+aDr
t4ot5jmsZu3EpJ1k7UVT5b2sXk9ouKTfgfaA90q5oXzSgB8gMftlNIiLMLQCBKjL+GiVBxhhLGwt
R5WwbM29rJIRDNh38WvhjV7g6mzp4qdW/HYgEQEcDwUmHezuDZEKj+nM8/E2LdpQkvoCAmV/lNZN
GJDrWZvNsVTSM2s4CiCsY6wqRFuCLkVxO+dZJ2KatShS6l8JOM9WJW0kb4oTlM8SAYlxsZPUetWk
nzP4koyRiIJl8rCKuMthZVHD4Yvi7jux4r5cfLivdjItKfehx8opaQLOq4MoHuvkekKG7wOUeHJH
/uE58BMIQb0e+1CWT8XuHX7zeJE7GaexxOdk2mVkOOssmS/ycWzlEbVQOFqDjUxujZpJOzODhb0s
dUAy/dvV4Wahq67c6e6xEyrWk89V1Sb/+jX1b7BgqIO7Su3mBD534ubtxxjCnc1VPp5Av7gfgVhr
Q9T02eCty+MSZ/Lqe8trTxDfuedDcX1QP/0wK3MB2TnsRc7LI/1N74XCK9TARh4yn3N93FFfzc1x
4xHvBBzUdBOf/9YUJhCVT/2vLqPL+3EhT0LnfyQoKRw+ELrVSDLZ4mxXk98UHm6qylRSulCTHVXr
XbhwhQwGTUTUvk1YN1wLULmlUWeGsIC/zxsMuFADDOCwe/yN2zmkRfu/ITrVdmj+Lk9TCzND263t
mHy9dmvQ1ixBbCOpgf0xwL6QM/Br+EqUBUwZyRS7TO2UwLAviE5vH+GBIIVCnNb0u8chfgrhnTaZ
r/12pvFpD43IJGrJcnxDGDE8hyAoiG3zBd6GcawUdG5ru/xYepKvuf17DVywgWn3THf3ax2tu1ga
4w3yQLHfJMJ7j59NC2jiBqQ1nbnumFcqYnW/NE5T5Dha0GNzS866p/XHwAZTMm+8exgZChwwvMrt
GQGNvTi2pLm0W6WUGo7u1C/vqoBKt3Ij3quVYJK9IPJ3j4Rx4nlaJ5IBl9TXoz28RwS2QVeEqHPR
3Pj3Z/hGJ6oHTzIYAdtlQU3OJV7p+Ug/U2dAEDSKsULhdjqe5PHTX+xKYdh/LSqDj5tclZRlZoqs
3NTM/mNL6+WXRnkXZTmIxXlzMM2Mlw+fCtJrAkUVg7JP6mTCHVBC/zNH+FjjoPwekinF2WxbpKeb
3yY6KlS8hHEsxeYFwk2SN0lLzdh9qbqcGd9du+pHXzOkVbHboVpcro4ehl16UoK8Drsdb/KmEM4Y
GSi6/uRvmPzC1yZmEJ7anmofS/qM1N/H9ptAZKALBlRhgsxcOp7G97y8079DmkskRXNii0sQ+VX3
zels/aR761PUobbk+c/oFUMkVb4aX5ktLjbAbmBuhqAUKYz/0yiF7PBG5uWIpLBgsCxmznGlC7bt
Hqc37dqiMxz6tuqV9wABToHszSK4aVsgtoh45ho0Mt/MU6yvQv54RWsES3FmMBxY8EolSs1BDbZl
mLTe0l+zBL7I7ku1xPBWqqiCQoYZzvwEtSn7zcJ7c1QR1J7xp+QwoFRISiCoPhw6SzbkXHPwsJqZ
Scg7cxi1Jbjsk/GQgvn5qrScPqwiMmcTmgBukfU22/llXHWpTKjAN5rXYS91y4A2KbzeK+2OpTLb
6iUR12zjkJXqN1Lw43vxSsGdfSZIMzJZ9955Vrga185b9OAJRP7G1QqoOzlo6T6u23nEq2FM7DUS
dsyh6zsnGUPjOirQ1acXbB0ydlXm+FHAtPoxOFcB04nnD864KgMVu+22NAClLow/DwFF/+CuyiJT
6IBQMpoNYxjTIbmVsIPp17AjfqSvd7Svx4AdB+xsySI3mEHbYf01XS0k4Oe9DFhoyxW4SveoXJpJ
GT27OLOTxhayJM3FCIr/bVfyh4WokGNjEX8tCm9JVgl6WywkDroB8LNZuGaXbepJVDZKO4sXpo0H
ELRlBnGt2UwO04QsQI/KEL7uzdd1qR7ViXyOSbrGgUFAgWZdydj7MH78Is4QGw6YwRwZkFkHofV9
/VDk2Fxu6QHLGjh+kXCYo7IDitF5M0ajdsbRs39n1mP6SZJsvRgvbpfcynaQJOzs96vyEr9/qtuG
DUfu3DQ5tPpTfpo0XsDiDMjgMwkzLHkqczmyLrK4+S3mAn/P14pRCL6Hhg6B8eiMCp5C1zE9qbqM
5mFWLw8AhjdirwZNAjqFPa6xPQOj3YYN+ZjH4KwAFKt+3xAntSjAhNiGD0l1mFjDK8ZPQiXiGCrv
HHJIYCMeZrL8Ylid5QpBsrpuBlbEyiW8MnLte9C8mB5DYRkc5FAgvOeSSQ35l9qfqqQIoEjT2GrE
be/5mvInJvivCyWykeqkp/G39/+olzRSMgOCc6bGb9eBHqtE/PhUGplYmMz+aOlxJhm/mXHQT+XE
EAqxG2xZupmr7I0l6jMhbXon08x90+iPQrmYC38IQItDLGwf2sWpDa7HuO41OVRBmyTrAXTUFUX5
6De/7iGeW6NDvUlfKjqv/7Fz559TjvjqsI0CPwTJ8lEnpUuEouTvm6BmxC8mAlVGNKwQJ4GkYyuj
yHSzodFHSXVHHNVd3R/VxP1Sz2SOjWey6p9epTT9tmHl/AUGSbcj8IdY0Vb2fM0jrSrYhb4KJsbb
7mxyrrY1CqMDuLDwvXbhbytiko/JxsmAzmmQN5kVkWH9Zyj8j1CEbyVl7pKqFKCfbrF056TNlyPi
fgWMZK0vy8wbXFetELI8WEXQBfCQzyZMJ3zsGIOd7wupRJD8Npn7vu05BkNsGWJqOcES/yGrcrPD
wsQi0K+6agSUJ6fWq3wVpDmEXDKmYGMYF1KdBL0UDDOde/fZ/okGgG0na3L1TKLNw9j5atNFiTpf
DlRUyL+3k3Jno1ZoxKB7WcbUAvFuV/dyqKZadi37zteL67qONyBABOPLYwxzgLm0p++eZLW/v4OL
5gZvAfiPGyJ9GUcEstSXT8klrj6Zumx6+oSgUiXT5OdUx1wkAnTexF2BLhXfAfklsZB9zOO2ERik
NcrciHtWBag1FvsBULtsAPzq1lO1S9mGY7mLRaxG6zTqyqJ1Y4P7OZHfeqoa+SHXO79S62Ary+bk
LW8e/TRha/I20Xa1kEGpP6gTftZEV+SXPIz2EY18JkyEyJqQgysaueB7LRaWL/1dsM4MWB8O0MA3
xpOD58WbsIMlVmps/J8sJWr0bCKIueW9HVJel6sGE/K5CrtBnYH6UfsahpgRzHoVIPZM2jbQd3Yd
bJbd3FryQTgiDAI/iU7fuZXSMmJ87t2reNSXq/4PzglBNVCSKKZCI7+57cvFFOT1bsUp5PG7FKP7
r6nLU8D1xQfPsqxLEexGJOrM5G884E15iBoP2+hdxzBZCNCgBsRJwFQhN/ZiswSNgVb4leouDBeo
xSbJlVwGW7VZu0wt+FfMZ9qG7phHUs1SQ6xMp7sNa9mOfTAlxDzT0oCNl52B4Yqezkz67nIJwX5J
9UO2GqySPD5E8ATYvY8P35lPVe3so/KOCg8o6F4P+2D71zLjqzMdhCY/AKKdlLl1vVxQycrBmuGK
mI3CxdzDIdqMT+4ZDxI/zd6F7jL9pPdDU2vKZeChTpXjIzLqy7hVcGDzSMxilCOEZYy/gsoclzcl
u1owjqAt0xIkYFulgQLbUwsukKsmp5td7R30FGAvy5YawWTDA+koNAfja3e4ZyqfhFHj3tkVnp+D
JqkMyO4UsMdhaMPSkYmlrsL81uZJH7eA0t/6CYKc4v/iGNnT/DePXr2ik0uxAx/7jL/5CdyJvNOx
g+8sMlkf/Z//aKjqRPOPIjWmo58GURSR0uxJcvSchiw56gOitPE8Shkexg1UqbaxnK1fMmKSOmwr
BQmVSuxty52Dnw2cjbnnLWTicb7RtHV2JhlaW012CNVUKLVgCd61FFNa3YOr9nWvGIltoBMEjJOI
WfJDImuhpVtPNfWkVj6ueRi0Svjws9M3VDQfkI3gn/MvYOwZksBiSPqoZ2YLLObni0OAsjQnoGlZ
zXbC0mgg4FXiDqE8Hc8Ds39O6Ygn71FAuW/UUOmOqEEnlMS6a8gBgN5Jg2rjrMS/GGJC5/7kFV00
qQT4dBs1LTp7AqbctT6ZHXVgT4gkFDHBbSRmUyOTLbxEh9Mxl/GKHTIGchAImXzBe/QtK0LvIHfZ
Gl8rSgnukStWwZ4K5BRGup2rU/oNFMQnByRKOVrqVPUqyiZhDJ4DIGx8qdKB23XqDHnsQZmmQyQV
a9HV9qdXjxD+meJbTr3bw+Z0G7IAIHlidDOEUhHk8FuI0cUjz93AhVQTJthQa1UveooDDYoMHlUC
1qWd1hAT7c4Cz2WHdnXEdQKHNk9pBa+XWLKf1aotrr6UMGXYEUvcdNRVuhI+RwZw/Tn8lkfUMp03
DNhMBY9I/+f/Sn72sxal63+EOl+8ilR5Pf3jiEWWrjWROK61RuA2gZEXaO8FyH/mqk0x6DmVK62h
eJ7IAxKaylQYKNNgtQTypQABc55ihsuSh/Fz4WZ7vCSPVzQDeebClHlSS7fVmqEIPTwf7oEZGdHh
kpfT9SKoyESwe4xlVCk2ddVzxnrZ+pYypewkzUGwRSqU070WTDgcseA6kO2V0KtMq7VaR/GZiuo/
WPCBfTTbQnjSS4GeX0AukJtPIhqI7vJS7y+W/HPY8RkvP8ZB0eLItp5eMMFvIow1ng4gxuVLFdOz
8LTG2WtCAnbEhudtk8fpsEPgaSdwbmn6iVctVzhfeWF36/RaKBahtjbXUT6OV4MRzmmVyu/KiXIp
h0WWA2oMCTnf007AwxQ+dzs4arqiNj9HK/PrgoVfYRyiIv5j5eO21AuZK1uqK2yqw5ffWyDrc1Dw
ZGPy1cw+RdcLcJrdgmpcwQ21JrrS/Sm5U2gLIKN2i4psiOYIt8sNjvHhBrS4228qCn9WibsBsxb0
anbU7M49cdS47zq4nAM3AB/qvULtTHlR0+Y1fj/ErMh1Sd5/8qXihGg+E+SncSPujn4f5n3j94Pd
jaUuOHfaOh4QUV4p6GXogpMapJQVrHZ9FLUUfbCmIn+Zz+v1dJFZj71jjTukZqRV1PsKwncY0+Zd
5DoDZ81EBAOUVLvxW/Awwb/cl5xOWdUxFMxyVhLzDWY2LJ1Eo3tVYdFzLTz5vbAym1E6xBW+Boui
rIqAzPx1hCSSsQ148UBrq2QWGYqlr4EAvGBEeTCkAPaFwLqcE21nUbI6jwv4teIVyXELcYjX0YrV
fueOFN4sqWp3e/lEh7cXt8AQJ0zKcaBhwJmJC6ol1vNy+eUMwQ6fN1hBaxgCn1ad16pzFhdqYnMP
7MhF6p5avl6/7pDHA1uRx/xEwnsBYfffJRxNAV6pI2fJpmvS+rcy6zNL9mJka+2AI7PwUZhVB2dZ
uyEbbwnIdeS8p4fTVpvBYRobRxlUKokZCbK7U8A6KYYvnXbUJA41Xx3dXQVNrrPChotJUNEmhYEJ
zsvVhFO1AKxIzoogt5+I9uCvF/mlt8OPm8AGhCoVhJXLZEYNAV5MWZY7/W6rqLm2P81yAmIOtDeM
BEYQ+tz7ZO60xZg2pOiyN4zKOohAeF2jCsb6h8fTtr+uVkxOQDiW5N4iIg0+xHx81lGBrU/JAKtw
epcKyhoPvKuOBzgYeIUmeeWvzy9lBnWGs2BFCL88g4GInq50AsmPvIP7WoPhD4nwGdfmvBMHGTmE
SKd3ovDXvVEPMWL99Cwc4kMOnEgkW3WJdCpQ+/WMmDV7z+9Degikkog90AZYT5G7UmBTPJc8AuFE
RaLi2CubOG+D9hLB4WQ8XQ1DkfPhk3AmHEDNHcRaybV7lHM3hMkltzKkM+FgqaSvB9zm9TzniVqc
kfV52EcWTZJiuRQ6imKOBZiJ0Bgel/MBUhEpyZQUgmlOo99GF5n/zcbx5ki4yNieaPea4bY65U/d
BYWumf5VilF7TX2jWh9Zr4tq9d8iuI4Tdt/GoZDom4dVQFswGyuqSxpj+RvsRQl8ASj/IzWw/Vjb
q+X+rmyidm+IVvFXESKwAUUkZoVx/H1CzF1L+RnMcHXw4tKJ4a1Rhf3SoiNkZq4wX+XvCULzs2Ic
A3SpkmC5OAmZe78FlryiWbJJ28md6D5/nFnpiXwx3HZoREBLz/a+M0J3RmWuwmuvu56twbVRFys/
TWxnUinzb6tyMhfVl+eifzkWonunthRaFywcFd4xbil2tY3AIi71SPeZf9zrrH9ZRIZ3lJEzG9tx
fkEoq87e3BhqKIE7r/RYwxbyQYuqPP/WKIs8sZVesYGynT9tmina0v4JMS0DX/6zAhxrVq8y7uvI
PY2rdr1HT0SvGgvdN4fiF8LTqZvS5JzF+RZQogPZH8fnhzlz/5A43+b/wMTWcU0wpoq/ySyZx8uX
7tIoSVv04rlOTUkE3ruWbtuECghhoFwV7xK4q8ZYCbRK2l8tZPorLNWmD5eNubN/AYC1tiF2ZXxM
B0brHQUANBphqIwAJ9sGd4H7xXqZMzhNscImO4Sg5Kd6IGu6vvPniqOe1jaxl6LVr4/pwiQnNw0q
sfBZnpXMBabdMdl0ifxcPujd1XinEC2iCl8pZs+dVOi+6nKDHJIodq6Y/NL/UssVWsft5ZGQOfpA
Gm9VjPMVrxZxzJF8rMNFPl3jd/nTMJbPpe86rKb/tGA9F3hA2rEccQdqexQqRmLxwLm9Vopj0nS0
5gMMHjzBIelD20IZ/CNJ8Gmx7wXNo7BcwPidiNkjBr/bRQIU3Rrsk3DeoVcSONdcp933lH4ZVE2/
x/E+ylYQ8cnSSqhN3uVY+hhA/QyWEnCoRsviDiBKinJP0/Z7W9zPl5lvbL4tdtVos8HGRngUHu6A
ewvmzvM6djnz10FSuip8xg4phbgsoH2FwocpE/ggLRlqFrRYvBmXUuB0vvL/PLNXpTtPGlJcBxt3
jwgRseL72Bt7zqxsQT9QjVeH2X+ZjYqKGH6IRnbGUHx67ApnoudHj/R67xp/rjuM8RS3YQVvo26d
4Nq92bSZWP/njviYWhuUmXTr5e8SLiUcYiMxSKt6HTXrWAFeVw8nBsQs347/CTUGUmptFrJ/ApFj
drxkgej0bDJgRJWePy6y/BhqwJ9crY0BGA3wjji7CiP/Pvbmx+gvWWiFYkO2bp8TPGqzx+N4IixX
V5JLPw620uQP+USDvbMv8o9dZfEjhWGaQx1SOO7wKcnj56HGTVGYfV0+e3qDBU6sKk57sTlIyD43
W9yHWZ7VpyjMrT7KAcjhGt/T6P+UUVCNvA19X7I1x4PshDpPEFJEvnBC7wy5qoJlqewch7pKUVbg
sD8zLcOQot1KUQgFNxfcmgHJc0bxwzZjddsTl9aqhm5Rb1c419K52/GcnCZucfqRK0/SGp6L5YKi
AXQCalWggpKT6iyAa+dg4JZKjlTEazYGQqiWU0RxkYaJUcodOnFtnqguAgAa7adnx5kdqmyIebRT
cL1qcn38kKAoxFMyDPVXCVGxLzCwEsSAXwY3oj0pkuov3rJS0lWf29O9aKT3+zCHKFSqsJAD9uYt
Urf6I7tCzqQciTuCLJY7cGxt0QXuppAznhAIEOv8EnUkG0Jc10btZDFcTedW/kTx3k5YPyaduiaW
Mpqw8qpQwQ+a0+JhyK1m8JJKCA/E84+rqHRyXfzBGoBOAqKtqFhwiUwze39hN5JyGISSZfMJbPPB
0dl2XI7PB2d02iTKzjSek0pEPXd9CiF8yfWs3UCtWhgjVCL4aBywRoERQbKaCk2SecoXvxsq3ecd
Rj/nZu1qw+h08hytTF3JnQemMCxD7JtyCVhYLBWS2fTtQ7k7WVpEWtNIjX/80sMdP96FxdZ2NSKb
BJxTFrB4Y/Dav2yb/QVpl0Hz+zn7bI84gA4x5UmpNut5K4QCMoG8j/oCEJn3WOasQBn1/F/8MPzt
SyoRKTcdLEhT9H6TBWzwYHCdFkx7zNKYQ1NFM9yWmda53DRieTzfgNL15N9SUsXBuDR671pxx7ck
uBKT0U/+CvmcSDkT2jlgIfid8592aXPaDy3X3y8BBC8Ent0g/aYBj82MpQN33P33RAvO30ejTyEZ
lvuLn03bzfZwLOI65UzWs+h0/5LyYMkOwt+9v318ne8DL2kmvLrQpktqk25+2yEUOFHdhWtAmUaO
/dYpM2K9LNNTY1GTNKm9icTE+cHIeLz09muJSf6KRDB1YQyh/W5G0Tlu167U64Ldh9LZF6H77Y5n
2ZLjnDt01j3eJc+vHJQaG4tNqg8m6XW9lNecsrGNQ6pIQVsBbqLsixUWZ28PnR1+pncuie5Iz9vF
XsKhU+U8jsnDD1ZjdmJMdgVhIDbm8cacE8Jcx2M5TmedPi8c5zBNHqffUmvgGGHVqmKOB3P2lMJz
Awb1gHhOUd1A/mIuVdDdSdH6BkyJfobyz9BJ3O1Y5uMN9BRE/ELD1I6oaAu33ihyaY0g+7/Cq+AM
o+J0R3HpXA5p3BblvodMoOdBQCj//LbhgeVovmEnzO2qQZauJxXNB5yMvVE5ZzP3ScbhIJ7V7XET
ZQabQktr/cglFJyREx1atqOTX7QHwVjY7Cht6hhUJfH5+08BuAZmzgP0oda2no5LjOvMoLZFToiC
A9kLiseDlN/KRfvSrQQE00mRnaYzM0UP4QSp0GNzrdwcUXF121FmeEt3LWGm76N/qYDsbHZZ6bzn
Yg/v7hz5D6NNz9r6UD2eZ3r/X2dfiSaU2u1V6m7aCpNsTjGVYEI3Yd9AbwHxG1+4SJinYheAZnJo
RZg/rIuCu6ucEaTR99LUepOuH0h2Bt0jgcwMn19j7qmVnWtWqRAnwTvaotJ7FP4yynUb7PCUPl/1
rHujrQxfm3BKWJKHHynenXaWiQDhbthlwXiL0nnPlL4AGrGW7RsADz8QiuMPJwbgtCKADMT5dCXa
hRX2IgZBNOpIvdfUsNFKm8VcvzGbXCU0HPVDqZfpaBHOmYGG8xkgy8zS2VYhoiGdAua0JoidDqf1
7jgvZ0GyfrsS9NIMw+yEHe/U3+V+GuCCtwC8WU/rlWy/S1f14Qvoxvvpg0SS2uFkjhPaEOZGDkjY
XhZWMJBRIqTgrJVmybOdhXXHVQM0bsyOYpzjhg9evT1iJygu0UdepIWq5v4W7/KZ4QRUtQnRNkcQ
nrVuAytOv8zBjz5Z0mz4hc16B0DQDjVOyrrPkvAW6oxSGKXDZ3TAD6VYXCTJNsjTIbxjqYdZu3Lw
R4xjJKK9j2bcZqWm8ZzKinZ0P0nj+pvPK8PkJOqZ1GnAqjYCo0P64qTGgclkfRSYZ3QG4Ye8rgAQ
norSQwreHEK8xs+uZy3xR+oRIzkMi2/2v0yga7hJV4y7UUpzRrivqHiKD0KbFbUpszUWaSg8E4xe
5vSFnxNM87s+SgtBkfX1jGMVQ+AiSJtpkM/Qj8SYnG+oK+L35fPRH/Y+dgrfkBDCQilf6v3+0Dvo
qMf2T/5TraZlvDnZgSR9WEESks3KVh1B/zpYuHtfGTHQTNOQ/xGitnr2Vhkzw23ix+3uPSJqiTiG
25XiGxuu0ObEBXB5WukA2t84y4L4AQu8JhURse8IQZiYzn4zUIOCVsDK8N6CpWk0v5dqRmzToPj7
8hU2nSryz1uoSAq+vhsvfXmKOKt0WLucCjtgeBIOHNUKF7ThrIXGCDDzkFO7z4+DHrfAqGpEbkMh
+eFc4L3nay6KhH09C0ONO7EPBPk80xVBUAR6V8VbaEs3ruzt1n/MSrqWwX0n8ZFkyKFjPi//6oMI
9glUOw1nmRTRDKgTyxaum2qkgsEfOzOXQC8ekZwLT7c/oHknreNITPrd2NrAGUyPTSvW2a2meNed
WB4cadXjjZukbwZKiJBpwx/hmQHCCu/grLlRKywFcbznB7TVT0KD89PmdVWs9+eCyFFq5wxu2R+Z
/XUlyAJnvGB3gHeBFAxDXUuwGAn9NNBac12bf/UvfZ1Zc0alZn2XmGksT3AKhD7mN7ci16ZWny3y
Gpmn1r0VfDL5hLC0TI16BUD8Oqyw6hd7zwRcszslC+oq/uBSGD4SxGFqGhC/LmganY6vlF1KmEvr
I2GmmHDi8USoRaii4vUCaxXbTLBJGK0GJyJhMjELlmAuyhfbqUVv7UezejjjyBZwyjVC7C+2CFlI
bf4l6RaDTDHCUes02w5c8Uip64VOTo6V4dKHvHSlVgONbZ3sQbQpwDvsvktOT3g19wKGn+v3u5ay
bAV4PHhIOIgcH2o3jo6aYVoj1oKnMPFKM2CzJSGvFrGPO98a09GwknRRaFQq6toThUeLydGHI95c
wRGcmKslc6Ocsc3CcrUsTVS2n4/k4JIhilxO9VixikHwFVesmbX9LobjtlbSJhQ2mbvke9yP5+Da
JsTVxIiOKyGwKxJER55BBebKSJ9A2VjCW9wCnsEEQ0PApQ33vC6lU+6YzItoxb3cXw/e7jx1GnCK
bDcbgH/gYYEIQTqGjsmmFKI70fjzfRuYAW4SqSt8XUobnU6Kp5TD50cPzqGpIW71PvNfI2sOx33m
Pvpu2/tfuslPg60maQbZCpe2L3fQiXmMsoCZbSJWWe5ODkfUUleDSN2GdXBWDabcmP8ENLhp+Vhq
2QqeRufHBK6dtA8uvMtssnPRTCNatv96wXuvnIhSXhvueThxyJ6PYcLYD5Vv7Tv5nC+hNKS7jD/P
Z+W9Q1u9fenivUwEqC8TcDkkqvIwRLP25xYOw5ZxKKMJirHFilqHO0m/ipi1RFANLQbBxvyFfbAu
w4BQSsUfSlpeUu4NSgoFNflpZFK6FwUnYjvHmHfiGc4hXWUdlRSrpPNmegkhQNqzZT0PeXXO4aR6
gWYoOnD93Jnd2Q2+WRL5Sg38dYVzWGvkwZvyndusZw7F07PQRfBkHBmNxu0fncPJ+b8FhApVGwg9
55OepsglRGaMkk/S25cXfzzM+8hwX1LxH7KbXklvJtukHBNreoTOFRB/nE1V7l/q9DRinjUhlBJY
XXN6H3F/Eb9BX84cspVmaOQ0rWoMIPC1mGrKmmfR1YDW+ZE2Pel5LIi9wR3HI+AFLlHF+QGwQk8h
aFR1KM09vPV1IEzumlti5Ka3yw7SkgUQoxlI7T5zMgUtH8PxSHPMBxuUHvMbOKmckg6qaN4rHpFq
qoLxThJvSlB4T1vjl/IZBnsHBqO3amFhlI0PK1ayjKTJnpV2tVdkAzqvWili5TsloIUbrOlU/cP0
qxE7EfA2bEoGWTP84tjt8gTiy9w6YUB0jnu7YLmECG8YNgRrDdTcVTP2G4qLYZC7DSZoXhn2nit5
XO4y77fOOm67n8QTAUm50QXOv0VD68Skkr5nhycpDZJVoaxg0Qa/zsJjnf6Q7jsujHsw+V/N0zhk
OnOyInj3uh+MUzQSgcg8g982C+w7F9Okkpp+a0zDxfo81yqviGIUD2pjF3OHAZQnMPk/YdfnCnzy
zB5szdmm83AqgeyK+UEAOhA+SLrmw4kZ7TJjcOPnxqd0PGrU5HPxbp+q+FdMMX4kYcyneiJp7Xao
Yv5fj+/Aj/epy96Py2iHG2fUhLr1/x9HgfJ04M05HazyEXNfBWg/uHHZZyHGG9rXf7W+yF3G+QSt
1Aflas0e2Y5Iay4T86X8/NJtCZ7cVcsriSYOnx+OoB5V8JSTJzhjzKimUpsoewyyvluL9/lTHeNT
rK/PN7BzkKFhhhE3VljAuKxgVTtcDe274mYM3y43aHrbSFkxACciTF8ZiALvxUUW9fYODL0dfHTY
t5ukeY9lpbr0+m9WL/23amR8PQvzEisKD+mRmEaJTAMPT4cIcIRIWugRX9iF8C3skBGXcSepOktR
ph0uDMRGdciI6xxBCzAMlLLavyYQXGLReZ/DS6pTZV9uN5WmkXeCzg5OB7tfRiZiLgjV6JTy35xN
N9+3lm9vUfNm9NG6EYlZEd2k56YNeaCxpLQ23SYrqn/NTEYFZJple24faNw4xraBY4mPNS4nAol4
rHsY9oFSmX04snm3lYRtV034gIScxKoIWQbGUl/LbAeh6/bxarJkeogJ8c/a2a5egODSKMBPWKiw
qv5nYKMs3Xn4Kv1q5Bc4aYV/4qzKKczGHexGZa4etnvqhtZoZEamNY+kfUUFUoTLBG6J0KRagsd9
6/e2z72xjrms5pYPjj/dRnFYl9gEs4ahDtK6FrbORnmvybVZyj40IeGAnUeO+kgv3yQyBiz2z4kz
5w79r7yickQMbHJOQ30Z7Ww6ZoFHKcCwNT00Y7waFPMTSMgQE37hoHy9JnvIjgOqZJqcZ4Ylb+Ag
g/y9lVEJKL7p72LbPIvj1us2ir7G7HucBnCk80hM0J8KcOlHZGzmDi938fM3ml0TVJfM5I+CXK01
Iw6BVeUtlYpj3QTnFwksFQM28TQaemZSUwM3vVnp+vAa1s3eSrr6J5rDUHm6dJ59LFmYgrDHa6Ny
gjNqPxV6aVX528JEpa0rfAX39MvajQAPvwsP24NwdCZzElTez+smbkngJygn6xnCdy9OfWpFKpdR
GRVbBUGiiuppXIPAE8nqAf/nthAyHXSRLNykjzDq2kKO9F/L/+RAIPZvobeOhQJqllv2UydSyqL7
7eqCjhrCHNLmK2Y1UolmWLkO1gBskkpplGrotRFvQ71UjvyYEbvpA5Z7SYUdx3jgfOM6ymyPRu83
zY+CmVzc/sWTl3y6A2veKt85nsQ+3BtquZDITjLqMu1gFB8nPrT29QhGRwdsYSwDoXY0nZOdabrF
ZSUVt4r/8BGZV76j4u9/vsqV2UWVuAajlLOglA+jTVPaHuOvS19kFznjlmQrIddxSxN8jd/36vj/
1QKuUGuTWsKzWJGs5Znmz2rJLMPcTKIq2SvQUXMJLP4zA0476SbUqaFAiyT/wbINRbvfGsDerfRs
NqpcX1YZSCqJlF0JzNPJ2ibRAnvh7r+fu9w1NlYycFfptNd//e58DIzQFdspRI1IaEjh72/G3ooE
QabDKC73SUZVHXkX8XnSAoBXAM+q7rh00dnr/V9yk2ONGCmCduvWZ/yZwFrwRjGYbE7C2ZtWGHuF
Xj/uOhkb0l7pacdHaumzV1XEOhueM2ta3iBskk9NdMkMA43r8MMk0Md6tDKHhfYCmA6Qy4b1z78/
70FpXdKBlw5p6yudR6hISyHhqJWdcmw5t6e1zjw7+OSiFW1QgQi/Fo9tvTvhP406YigHIjov7S/e
wOSASongEdzsdSLXWZUKmKh7Qnc2FkIbB3M2TdsslojOFPoCqtDKuU0Owlzkt6DejHG1TEJAsQOv
ty/G8DUBeG74Wi8ALRjFv0yQpxm4wxy6aLL+ciX04mmkGYkLxURXfGtLoi9RrRtGsDsmVz0d4wW7
TZleowV7d+9J7J6S48yqy27dXsOhkel5O79bpgrdjrfwMZAQXhKpT2+ntkaGBp+mIYnNURrRbiT5
GkbkQWK76gHabYkKPCVv6+2e1azqpfs9xDVM/7p8KYH7+6ZMA8f4MR7UDVEnls+Hta2TvFRkwc90
kFsacTGobuF2j2qsFzuiitA+or2xUAbv4yay+KT437k+ItC0AVzjUfNWqW+QVqgErv+SQP2jQfvn
JCA3KiswWNSDRnvsC8YzeGCZ/6fwJ/EraX7lK0bK4R8MR/iKyhYVSMQKw5gxgG8bwIVYA8L2F1Iv
IcG8v/kw0W8kM54vOp5xO0ZpUgODmwiLHqKPGsVpq4v5tIE4wMMELkOAjDBvFJ7z7aTHC4xVOVPB
mVLsq7ajGnQecg+f3tz9SD8lm9neavU4HeNl0d0y+Ts9/suwkzyt5p8FC5nCkrdnXacupfTlGDiK
nq6avJ97x/VlPrGgamudaEX9BUNfOpMyRJ3CmlsjcI/W6zlesXWPBgw4s2HMXy+Qv0X09Pe+iBGb
e/rLX8KtXxqZmAGX4s/FF/dwfMFxoP4epYjn3ntKmURIDmJbKDZr79tS0wVlE6hK+6GOpWqX3/2X
NnsncGAxFJQK3QIqWKIatS97bEkvcpxl3nsPvGeeSUSTLZGUmU9NG6m9vTubcs+mVFHuf/DrgUPM
VKn/P6jK9KqQiHLrGoEMzguo/ccBJwepiRd215LgkzGjrcsHPc/JOI+40WV2n4NirgRJJfN95kt8
RKCDSasciF1Ww+osNU/ViObm1T3DT+OhLNkb6H0nOHWcasOnSmdgm4nCCSFrxRoeA7kr3uHVQPo0
hxldwPcbVVIgO5bkjKQYje8QvvRe337plxXjCfNuEbbc75JfeTUJduz8fItL5x282gS0Madg26BZ
7PMoqHWRNllbkAtx+g9hDV0ngeOjoDf8FEYwgQvXm02rfXhuVMcSjUAwpf1cUwP4M6gHGh0yk/rG
+u9zwfxow1EqS4/ohpXtrNshAh4Jrou1x3WBEsFssdVZie4WG8MZ/kLEUsfka9FQDWeWhvlBdH3W
xR1fXGf4w67nl6DARjh+RqB41hjTpfVq1wsu9XldnDd0v8k9trcpte363IQSbmKxl6iPubOwCxVg
a+nuWn+PmyFxxYvyBdNSjI5v/PX5mtxPXuGOtVmT2PsWxcccYgwXz4nfvhtU1oLoYx+H2vf9W3C1
lmVufsJ1gMqSMHizRKuggsMGOGBvkCYFRtO2tg6Qvau7u6+CM6SUI6IXC5uIol1XW4N+3FgMxSwt
11SISexWaGjOiGO9OhknbsHNwtlD827iJrScWVs9qFVBGU5y4BduhLfbdUjHJx7G/YkWmevNy7bs
jS2wkJpi0kgmPVgQegqi1Vpjrkd2NUJ1yQplUcQt9pf7NA/p50uHQIIML9IgDEfLmgRxC4fKCUQs
9AQODsvUOcSL22OI6oS1wrdMs28OatTQOR16mL08IEZNGJ3V54QBuNfTEuppykZoNYavGiMFL82w
tSYowD1Bjxf/LJLDIZkSn9Iv3IEXQMBaSHw9+sXaXBmzgbCe6URSpsdBTUhsFTlvqT/KyQtJboV8
geMjPwAhsvEBDnFa1O2gCHRxDBdxU3pCFiWj7GVXCVIJuRwxQA6VdwqqUbM6oewVo0R3yjcohFKM
n0+UT67FquMyLsiwt4qExwiJtlPBW/ZAq82K1CEOvksU+h7DJHrORZvXSruftlVbUUwr8TrI2NfD
kImd24SkHxKfkfcQx4VMX4I/BP9iYdlako95Dc/u9t0isR2yuBOnMkUvf003JSyd6o4Amw5wxEOB
IU06z4Yt24JE/C62ZmMgaQV/2bFt9Zw0KY7qmazFB/xLE/KpPH2nYgHo6RY6BuA3qLrlMm+hHwyL
Hck8OuKMqo+gCy+54xLPJHLOAvM/y0Tg18bfBNneWON/199lpSV5Ao/8snYlZ4fjYLJTYlgYjnd7
jN6TwAaFlZ4hUFgwTZeEPJpXG/MsfRVVjyyKkv0T8gSr3hTBhmPW443Mt+MDl/l4cILiDZvlZB5q
u4EsudU1S1P80/DYg9wihcyaZAuYRah05ojXS7jrLyGKeazpLv6SslpyoksKj/AyZlXkFWEe6uHn
F11FnvUnKXfoA+Js2hdF2hRl9qXuRRv/HgmuSPZjOpI76aze4MsRb5dNTQc4JnbY+Br1f4C67oeA
VlBHyn57Lr7VPmrQ1tVrVVC1veVbUvQg0NdibSjnlCsaw5RXyDHUm+hD7kgk/gG5qzcV03wjwNps
z5jWf8aHOlDtlTFnvJ8whe3Kslvs1sbMieSO5Z1Yi++Zqj0o9RW080+eCW10Ra+EdZj3RLWdMMQA
4cHJ4j23VKGL+JMl8HU29dRP5nvRTZgtFdmX57/6re/eSBFUG/Ez/KzxOM+6m1OIn2rOCMSY/Iqm
BYaAQHiuudXH86/gHmP9JwItSZMiQZvWNRMe4+bO5vB+4hl8jF9xIJ1DS3P2jw5h1Bq2GJIWhn1c
CjHSEg4V4o/3G2WReZmjzIYafwT7TN38El6PDGOIoWWz1jELxX3Qf/QqKR1LIlABxwEj7ctxPQod
3YLIvqGGJ7x4FFFeOACuDQRHxlJpIEnzp4oPIQ0q6k7fHWms45tZCXvx9HP6YIz8Z9uDt6W4e+qd
SVRexrwh/orh5YWv9XGd9snmWgmRgbXy13mtXAhAtCuwsQritBkZ9ncZaOTs13Lb1PjP4/vkQpEI
1VKp1YuukK7ePQtG7d0EGdG+q+8W4kxVZkK5LPES9ZTHGpu96S87x7qczJFI9HK73cRLjsBwyxR3
Pv0CRWDihL9vgUb2YwLW4OVms0DNSh+/EG0yzo3i49zQzvEkOrgnZ6MMF2v3PsV6Q3FI63K12cou
blwiYQSsPMKEmygIINl1GpJFA8lmMTONAuc4kSr7534sBlLhU6G0PypMVgQSff52H62fwmVQGXN5
u0cmoSThurfRZsiPfSwBSLnpQF2iCwxvDesAyXktbrZ1n+NjQWkWx3jUDK+dH/NzYoNL0nBe4MVh
lJi0lnGB0gRjbn0qn4W/4IXPk5Aw9uHi86PrdE/h2MzQ3wl0gXpSJ/S3NRqEH5GBiZucBh8+brR+
rnn+swIDKWorAKBOX6PJ91Yv7CVlr2rTXpUJPKbH2wfnRnck3BzdjG3nAZ9SmKTURV0KZhEB298R
d2XPOZdjnHPrZTKgIz0WQX3sdgkMwtxP+LqxGPAdwe8w2S+ca2GpRGS3xInYFrES4uKVFKYmbh8o
Petz6YvCMZ9kbkNV1F5QBflzxg3+cX6XXkVpmpO6MHss1VBtMKGRK5YbMomgOxXRC3rld5A1CUA0
8AopqKnay2OX2z1dF/ZN/ZecMOX2vWxiYJsw84FkOv2gTbLuNl28ns5dYoz8hHrDw1WcXPOpIWc0
715WRJ1Rchlju4dX224/gVOLU1y7nyTmgWFPh/tcrJFAdOVWRUD9c38p0xhMjrzEPncTTJ0ch4w9
AP/xLD7FXuqL66H1BPfyN0UoYbrigDKNM+GmSgvnLKe4BUfZm10rSGZ2cbtbBVvxYxIoV/fYtuQF
zK2S8Df7x2Njwb4V0LWiXWLFFU+Jwsqp8NRPp7bQKqrDgym9tGF8OpohPCgnARjFVTycpNbQ65VK
XqzGiUx5LDWhE3EBn/vIy2J8hcvRAsNNeFyh32Gv1kiUPHZ3cselN2sRyK2hxZw2YckWq0yRRHnZ
992y6WaSv6sKRr+Ie+Eh/RKryZSo8O4c8Wxw5tDts/jgXS5VhHRIrjg+M/eDHKp/Mm8GOYm0M/86
iTOj47pt8Omj+zqg2rlxv7HJY4Q42Gd53MZEnBAYMUR9rfqcFsVtfs/mos/Fr/HpcRbCGjjHYBlc
fFAen0l81Ql9YhMLKFj8klmaozynL+yOEsFU6lEI1/qHnLSQ2wcEEG1cLuAgVi/+eTz/6wZbnsFw
oBlYxwdo2An/irhjAWce2njvGaq+Xe12mjtpcUrIrw2htf5sKZjsRUPiyyJnFVzkZ2fEU85MI6de
ic7sXWO7arwLAmSOfoxJn0wrGjemALiBafZp2Pk6i2n/jiqS/KYACdJ/W9KfhymlPhN4R2BNZCWW
wOHibgnZS1Lq+2jPHKdMDWOk1+sEKUR0EubXUPSGMwG/QH6xUNDBB2tbWBgNQQZNcjptNasDD6Bs
Z+ts7WGDTStHooPSjjemlmJ1E9qP0VncRWPv2FIZAYH/xSZxSpKb/R3pzVHtc6JQ80iJBydPLhTz
PvdZNTIiV77RShVcetNBE2NLlVW3La3nIKA+FobojR3B2YQsPi9pPlk84hIa+SdNkepkhCXgUuwC
lFlN8AZ4wKVIINpn5hSYPOtA8LdkE9cMkOleFCePk4L0AjeQTI1bmLPBvIM6s9k4GoJ3QgP8ljk3
b1z3X0y2/4Wa5415hD76JX8w6c7AJadhzAMiiv1u8aSXzcamft5DMgcOHKNbJAKyiYTcdbIE+eQn
rPO9IXQ4URtc/X2tjaCbfP/m+ADt1CO0jdGVFEnEHwwmidqy6/L5l1rz7wyi34aZzNRnZ/Q/hpr7
c/2pT+3HxdysZIQuMYS058OAZvVhQJKDLJXndue1blS3JJ3HKs2xACZLACvYxtq2mRERae9rEgtg
2f0DIyBVNGJ0/e3mZ2iiiVn06VJloGmIQ/WpxP6fFWPqAapWwhUcCSopAu31zpxxrj5oiZAWYcC+
WvI+5WChZCf1FuvN5P0mje6PKvBWvMdFUij99jpiBZUMosJ+4ghreKSH/Y9Evccut8OE00EC/z2l
G/YE2Z7iIn2Hk2ZrntZAoyHdw9SNfrWl2b8INnQhux5pzFIuCSO0NhuuQKJvxcaReJVJJMqyEO0O
DiF3KR1s2PrqlCWUbIc4J9v7T+QO4HUbeLWy+sKkWzfIoC05FJAzuY2zEbeYZ+ESaUdgt42V4FdF
OwLdHJyShQd2z3OcExhvT6W5i5sizbdYGgNhjzrauqbJPCr77KyAmf9nczUSZXmrHLj9Xur3HmFa
trK4gyvPC5b7754cC+hz9NguI1k8TMaZw9c0YLofNSuzDa7W72dyPb4ll60tO+lFNyIZwJLYQyAh
GkZmOsreyxeo9J5GXjItV9Ju3xSB7EZjOzXaWXeBfyK6QOKvZQT6/wHk14JXzEgU9Du5GEBRkQVW
S+7Z+awXaFDC20FxfkHHRdLAHblTGyYZtp8bFchAP141/5KWSAWwPMIeDmt7ggFxiF8YkySjSF+N
cBIcbu9fWUT3E2dxmQ+FkDGAi3Ba2By8+X88+GHId4UEofD12lCy6jIQ23w3/DfMiDk32IyNoJfH
hW195l8TIm+3gVsLd5NSQJBOLWRZ2hkoZTA1xAJZQdLr+NxjBoYrGlEmIvYsk4BOJUsFSs+3OSt+
47c+x81wxiWfOnISusbqD/LhSzeFyQrWXdWS2uZZPI9+3yoSngEGwFK0BN2z66KpsMb0iaoM98+Z
xM6y23SkM4jTBwwrLriepgB9urBcV76BoQqpJvijm6EfQKo2cFf2KskBby5c1/fP+ydG2ArjNCGQ
qlpcTFenDLIBTv/tgCMd/ztXd+1ngUkSF9gmVW9mu7AJ/pfgF1Yt1T2hq6KIvyk+S9Llfxi47qHw
uKLsoEvLz8ETAwnN2FmICkGNqs26x3RnQM7r8SMGYiURmGGruK1RmCFJOn9AvmbkIk+6WxUQ2/V0
lXOLtinyjkLSwcI+6QMvSUgzvUjCt+IMFwTO9QF4vAgOzg3+dvU0banQ8pgfqLoV0kllXSZ6glFC
jqor9d0e71V1evAppbgBp+O73V9naqs0NILXUZA8NxPkG4CHLayRs9e7zFA8WKqUNXTnzcqBIXqM
LRb5qs1YcgKVyXigkfBvA36jnjywVGhTBrDoEROon7VX94QdfRcha5wXwc0+iLr1ovtleRZpGKFZ
ds0Y+u0GPYLlpcr1VVSdqq1qFZ6+BBXzcewo3fdoUTVZYp6jY57dz3CTBqhLckucSc7F2VLKBUM4
qoDibltDHYTEWVJFoupgX3YmLy0U7YwigPO79AMFng6bvjnyw4SblbwAt5al0WQibIL+3PawQ4V+
XvTzsx2Z4Dn7oRFWCCjUeYKlQtW+hkyVyfquiVaLhm/+D3k40UxO5jeao6gDlxQAUX0KTB26JtJH
pUyIuoJC1FcmD7LYNkg9zj2gsSLVNk20zeM3aUfZMd9hUnBYmyCOF/b2VU60GCZYwNsJMv14fuqG
F5+Z+hiB5XQH8D8Hp9rsRmAr5b6NklG5VmopxetaL/ZiHfZpFv5yho7T176zVzOLNjJ+oYs/jw4o
xovmO3GfmJKuPmVHgLZ3D4ubsm6xAa1b8rbUDjsyJW/GYKSpjmZEknkn5FBtkwCpwxItgu4RkfhU
N6pgi4GBSPQI47EeudZfGXnePaWjwxWWOT3BJWvvSPYHj+m6yjyAvmUlc6MnkmMG737Jb5kqQr9S
UwkaImSVeYtMxPZKHOmHIKbvkX0wd3aPreudT62W/Twzyl1wucKzydu3Ra1x95ONElUN1KTmL7cn
PU3v13ufmcw9okc3k5pZcZbrnuG8tR+YGhUeWBmKmIv7cYVqrGeqeEzzP3Ut2tv8golmKvJRQvz2
CyJAo/UcBejbOLMKVH9ISs+D0KYGoiI0+CzwUnsIOusd/IStRegCOn1Pf7ujTc6t9Od9CZpGMKQO
PFJgCTPfE1M+3xKrzOysrpqYVK+5LTyoY5LQYMTjIRK1CA4+hRIgTXpQiqcXykmsCOrDhX0qV3tO
uMdpyNYFyI//sj6AqmvtK3Zc90Q4hM1v5kVDtO8zT0ImAjmxXdBD3xUUuza1PsCd5M9STxlFy889
3AHlXnCtVQVt41L1q4Sfmb4asxRggQVxOE2PQ5rQ0fjwTXzvCvJcTiEVQPD2CAc0U71U//VXrT1g
C9u3YeRfMYKTDewYz2O/a1bBScZpSy30kHUB88TLBgQk7S++VWASCP0VUvRlF2yZ0MpLao81bUXo
ZeRlKoCzZj7N4y/phltb1b7IWurZShLVw91YTsjRB2ojaW5tOUl8CZ5se31bxTXzee/pX/+wmsLa
UVGQEOvssrVKjB8GR7vEOSvmRSbcJAq+SG2BG3saDZG6jZcQRvp4/Pz73lzay+y24ZVouzltKI0o
nyYGNgGchL1ayZ6RIFTi2aKOYqos9i2jgrtWi3lWyGCbdWlo3d2BcZLO/7vkiMa5Yp584j8SyQLE
rdjImj51aQ0phlPT4EAjsCVKOciHDYTAHwvtgHThjHf4eZ52RqGPXpbKPHNQBitGN6brqDlsWhsX
zDlzUxNo2fc07CyOn2WsDDxatS46tN1BIWN95kfzS/zn8E/RLfu1ttznUgz56gYQNcyRlgHy/v4P
+kNC7kwFAw1kyDxdVq/pu3n+sgLYWDGSnqI2E5PY3h1+AAprTMBRrNrM5d9FrDycHNMGTr06Q5E6
4L7y96rqIOLOOkC4IIcwRYwlh7tZK0lHkXp417B8I6cMIGcqzEalkc7p76EeMS65zRv4TJUJJREx
8vE44I+xhUBW/8ew/2pMnkHnet7bkdVeLRJ8xJW1FLURCg1PX6Xe8vAQd+GdBGlZLg/S0SEdd6bE
h4tET/u8QLJiAvATRsJy1V8yLsxeqx8goxr6G4Q4WtyL0mVfkoBvOy1WyFLx/+BzU71IeRq+8m+l
7FQggvVrfiKM1hKLU2/MjX1AM91LMj30SujdTYgQtWBBU74EWluM+OYp7DLq/BnJTkhk4guArirl
Irp5F+ESb8S8qmFiIRGGBnZgposBzp63QAFPfWnfT0UA/lVa9eMs04Tt8ZqTN/u/+FF7cRR5ylB3
dWICcIaqCZjlzas9z0HpzSv7D0uZi4p/kh4smaiiJZ0HYZAohgMh7MCy/BILCZY7bThQWYYPbEpj
mh6SdcK2vGJHlnF4+Ku4i0LWA4vR1CmJFpupT5bHSf08RcCBKl9f+lNcBY+xqRB/S+UJd1AJPSBJ
i3kzvVtGy4gOr7gAeDHxtkC8DFB/fSlWHLQNXePHRS197xMchJQuHqSnIRamEorCo2SxlI0oFYXW
Z+74rN24hbjLvKaH9FrcjfviXPl9Vvs/07NSQXFftuGWXDo6jsNx6/JV2l5s8OHOjT2vVgRUaqG3
+ngFjWwFcsveAz5PUVXG7VAsF4SaUkGPpd3lxTpTgomvH744+4WiBMwxJecLn1f23bv/3oSyuIs0
9/vRVkXB3gW0D8IlZlDA6cQyQsukz8tOv+OsGY7+NbY8HCUD9mEuDQG+xV1nms9sK1x+dQ8XezIe
o9K4MIMwl5B8R1HDn/C6vNaxK8sGgGg+dRxAUWmFm9duEFdzKE1HLabYyXkWIYnfAAlsk4cxAPc2
YBuCaU4eOkqNcnTMgcryFa2wkw2ym+tT/mW+Q+k/oMhXcbUbYOQytp9y2kjGEhNIu4Xo340bfurA
FFv7LjSlsgvBndigj3X3dJ6PToeRzJsxMfJXxphK4tzSM/+Euu7/40WuMVl8qJfHBrFYySYeqBFe
SKyLDrdxemMf+gwCjlwZRW1wE0b9vwnz+q7bLbXUDe+VnsxI2+B3jxDaMuSEal9A7dIWWaAdqGad
hFXnMnN/x3s65qX0Ta/eoaOP65P2qEe0AqecJr2pDkzXqroR5yAATacgKg1NKHXeARHAalH5LZz8
LBxldrVwugNWcq7fpl5CcwaaJ40O4RGxlwSXHpWz/riynHRg8mdQpYLgs1NCi3tyHdGFz/s7XBGz
ua3/z3PeFjK4B3VL8zGajKV/TsJfPAJEgPEr0AB/gOWMoIgdpUsGwS5QUqyBLJ/f3NaoF4TGkwt9
JShZkICBXMRn+AamtOafboBCg2/K0jTH3LOr5I5odukLfH3942vEF58/abzSbPvMxF/TMnIgRqoj
UJTjWWwAJbPqdnZm1KRzxBlnHjB5MPCJIYW9Dqu2lMIIFQfLF0jjNmwNA1AV0fDx8bYgpgm2WVCs
cLlY4SaabLq5O3mCt8HMRRXs1rWARJvINrvAPH46l8lH2Gvxd2Cy/Mww/HJTkjh5Yxafr6jX0q1z
R+Xb5kUYaSVSlUSuJOH1/z1vfebOeBFsUhjowzD27dPWQMHTxKvixm6z9X9dQ6x4hn7eIeV60btU
7BibTgH37ya9W9DMXOYOyZvGYAfDDwKJyBOu7n6UkFVlqg+S6SsfArAaEVpSrZ3zP85m8a9EO9/N
nuWbx635pTu6mKedcezvSQkkYAZqCtMISqwdP5h1jfS824BRtRdWJxMiOW2JMInnw9CkU2HueWfB
fGDGJB09pFb56AdzmQoarhkSD2BX4kfWCxGQ4pzJuD6fQ4PCKCBmPATj6hOEpvGSJ+3F48aioaGN
LFeSykn6V0AX82V30tr4HAE62GxLjJ3/9PEQq4gk776P8JCKPpKUMxxBwNd+6kWzZ6LssUAwqlIo
/HaubRZIWhEFFVX1m3tzUUvZvfv2IeH+wfxv4EJTtQv6hPNTU2LOUDKo9DVbJf+0EUW79YGEO7kb
dEN9qzGykORqyUwW6Jctppen+xsYyAHdWeiik858e2+5A7L+O1S8A+Vb2CDS9y4Mls9joJXRSeFA
6ulGzxfGO860TtLwlDZzcVYHLiMhGaZV/vm0CXnqtdRavohcm9wJ8RVzVXoKoW6L9tkusKnKAph+
LdDYuWGQkdF0EL4Afx0ZNA1zzn1ESh8sroGaWKDUFTLV3Eg3bX9rTi+4vetCC/1OMoEWMDiOKooQ
fcZUTWgCvhhO80ycVQleaUlipFzWvQwk/hLy9QPz4EP8VdttgEt4gxUT2izKzojQ964k1nj2JAWL
hlruUWVrGQ+1IsDNS5LMUQDzhbSFbbkQDaZLs88vbeJfWRu7WTlm7Vu/e4EIwg8Rlm/ukoa5xxIJ
uY4uEuZHmhk7291VxXHEHEptWG+rfHNKWaWpCojmTACEYdY0CJtNqDxTFgiWTBstykrGl5uRmWOu
S9YBLX9FTaj3Ig82E11pe9xpg1H3QXh8rGn3oUSJlO2jhQn8YUx59/DcFUIUDk1mVeeOrUW+glAg
4yqsZPFWj1A1mFQ//sf1a3dojQjkG3ZYPFP0hNn84A/OYSp020MFqwJbizpz94f0dw3z906YLyKM
WXlMn1PGzaAHc+AQGnDvlyVWmsDGzcylXifXVIVtdqQyzkihtt1Iw2fwt8yj5HBiaLjdAHm7WabO
VSW6J3pAd1n6qdUhwWbL8NmBle5UQv6GuiTSbLACiSdHmsZiC7GJH7f41Lqth/q/Y9I8sAPFmyZI
t9TGrgzcutOf9y+fqLuXMk+Hwe4j3UiA3aSE5Kjz6dA+SNJ0ptbbkgGARDsZ2wiqL7Pmh3oZEJav
7NpqJmGmeX4X6LvvY4KCrJMbGiOrHvUx0zK3x2khvVABnwenHD4LgrjjGolaw8sTy1sUA/smzOOn
TfOBZGhlGVbOjzqhcMA5XxD87FyZAmxWfw9tBJrxCAveGJ2774qO3M31K8EBikMYI7kz+zmWIOAk
qdCGKeZgTIFAD6WzCN4NpNz201xNJ7eNF7UtABd0IBy4CK47qNE6bq1FkwISa64nemI2bFSosrmS
P8oubEDqDaFQd2wvod/uGL0snJEQgrUh84HQlJAn0yRQU/E0pU5Q/xkHwnZjmKHpkICSd4G0gUXh
7HsFx3fBmE0PlFgoLp6mrjCo5mRavF6dPy9EIwHMhuYMu0taSfhF+Ir8fuwHYzR92zaJPwqNsT3J
gRMS4umkLitRbKguOxYQdiN8DHgjdq/OPyBcmz/Z/iOggyU6NHNIi11SMHLggFD6exIco1Y5Ci0A
PkxIfmIHP7Iik5z+GCnHKJXwgSCqwx659fdqlmZe6KePmtrXqN6FYasPRW0Z4d7yeavTm/kjMfJy
w7zbBUaw1B+0HNkG1m+PKSCbeo77uO3eTi4g8KkAGWQsAesubpwnbF/Q2/qyqgb4NzGXGDvWjoGG
7xL70gATCFEDXYdodNvhnEwGAJe+MP8gMBtFpuO8ExbIrpfY1aR9L9Scrwb5vTZfmdXzAAfbtyFD
P1E2uLnpGzIBcMceZ6v0WcwQXl6Gkc9R2OR8LP6uGXcbD+OnFmjZ1W0sNFHWzf0JMw8iw/EZMQE0
IGI3VOHSIyfloensogyurQ5GYJ6HzMc17+CPMXAj2w5GoazEDm9+F00XBPrrYVxPHGilhqFHfMsv
prNg3npQE9hN/UCtlP3AztjZ7QMqium7PaNAnq6B7lOz1Rs4El/KSgqxT96QJfzWsPZJW3hNn945
RXuaFDf/1kMXA6pacgEWgV7p91ZRMYogPxyyCBZpNT5RrgjPNuB65B3HeRgPx4f0p8YiminZE4Uq
IM+IeTCQU9uih/+Bt44QMVmnmhUr3dhRLOWzBrHjoVRP2KGLxZDf6x8gM+BPubPUOe3/JLyPqSSG
orbEqF6PhX7Azg5gZlc9UBaZ88yv91Z59dj11G8TRCP5quw40U8k0jx/wc5uBdOlQe4Yjd3BpunJ
qpmzauwKSYNhf17Y3dbRpsj1A+Ac4GeV/BfNhV6Sju8Ftzb05UUlKN9uhFsun18AitMDdWUUxP8n
DQdTZPND7AaNM5Z1MbFMUSfuWtgr//kZXKrm5GDyArS1VpDxJE3NdisI1aWxhWzO/pHLcaWkGzYF
9Ez4f1WMpWznao0qK1B6KdSKUVXZBzWFBb+WMhj0n1Cn2VcErMv24l/jo9l8nLk79gr6ZKqAbzUE
Fxo6w/VboF5Lr9+DclDA8QkhciWoSI4dUsUvlsVCNEFLwDuhHNh0qQ9acn+Qxfqmvry6iicvZ7nt
z2u+qNPiGDpLBByklVqWFVKoBCx8ZbV4wfxHGrh8KOnEhH9c48vOJpiNYagoztE7KL9Oyg5/MMYV
VdaPCHzNe8sDSfNz5qoOnGG1EzS7h1CW9GimJg+nOnP4Qx96Qcv11LnFgAS/tMGqqo5zyX/+8LwS
QE58/FKcqO1tZT1DdJCehjgAsCkLJHXKifEAU7+JBxEl6PdMaMJ2zTEKJ/0lDH+yUOBAQiYM2vGq
4P0XGYMKZpCIfBXjr4cj/D0/Wzm1/TYixO6E39G3LU9lY8QYfjlWy3KYCovpACDefcOwjpCcQZVb
hfUEdKF+RSpCPJNunpC8Ah9PRAl2UC6l80enIgcusRvnBDdWB3T8Z8rhSLKcweYfk2L48KutlaL1
knGWv6BdzFPNesC8QRUGs+OSa7oXM0mt0vLhc5Lz1u/jf3WTztvgciQYekKEv3IybwOopBwhfLzK
ICxjyQrl//yryxFpDpuR67WU4wgHzMwWOEP+uj2BV8X9dJyu3qZUWo1rIDwPVLp4AqCjz7C6YMk8
6DgGhnJtTWUUGQaKhBETZCvm2StGhXHGAOhyPFWYDVVsrViYxkGw4PqL5iXakRVbuPnSMYX6IZuo
SlczFUUH5Y80BnVhrTQR72LHpbzvPMe3w+4NlCJKWfyYYfnHqxNhSvRcWVnKjI6OlxsgY5yBMiBV
W7+eVU9HLiE7IeX+W4gtyaUnAz07EA4NupTWlhXbQrw/u93c7NOCufZVrUqzFagNSH84erC27td8
nAseXGGVxrNgqMMsg9gWbBGViYAW/+ThrGjqvAkl6VqnVXgk57TlzneOz0T3jrp9f3yQ5ZuB+m8m
OXa2zKgUO8a+DbGvkb02K73RvzWqt8wZ3r2TRhNC3Xr4UeAEXjcqUyVTDCujZ5s6Gg0uoi4P/ZSv
UxSS/DSc1Wc2PIcnAMGR7efBHek69PMD6T54gmUnQ/Bvw6rcD1+umcApnViynP59GYLBxTalEvN+
ezfM63KVgG5Ob5sFd99WFyecTlAKfGpcgieqUDSqKEB3i1Rdz/2/x5WVM+jaZayu2OXl9q7cSb9l
upmCe7OBH0N5IOqMpWFROurHV3SDO8toNFSxVha09aAbODD0PkMJ0nZs77X/J9ntpz/3P1vcysxz
6C7EBwPiguhxUIuvoC6OgmUnkroaTzpGhFkwaEYVZnM64JM53HGZjYOqSIKkVT82pDdCUVx8DfKN
Y2iSBSceB3BL6oJsClhuKuk7t5Ke68GDN6rIo3+istW/5oeIVgeivLZRIPxPY0gFpFdRW/eQneIP
bHEhJTE2wEXfCuzhSXYSe7WAd+JoJCAtzLksIsKau0mpVUjTe3LYFXZykAhLSfQ58fYDNlCXFnLU
akq1nEkZdE19AosPMbEu4qBR3IGJw5DDvbyinH2O9KtGS+IlqM+EHaWBzh+YL+3Bjt3Rqmu6U5Wp
+B1iWfUcfVvlsPpp6DCxvf/F+WMxyQdulQIxk/lFjpNCvJX+I0aqCZDy2GdJbHvF8RSL2yMCSVEr
HvKXqZjfsSdV8d+lmK2sxYvc5osscGbbq3LAOS18hfp99WJUgA2t7L/YPSsIjnCT82wFAtIpsN2O
KBbW2yAUXwE59WU49gv5NntitEiqh7+ZMVk6xZOV2goP0LsrUs8v9kWjGokZ4a4/UZe9EY3+xst5
DosmECaw2sWa2F9dEokyHKybWL5GbdrO+3j4bJcHHCdF+DHmRgSAqZBt/Ztwn+L1Mu1Nrrl8keIa
yYWz9WnH63J+ZPcuj/FxH8FyBK0ypzguOBKIWF8Uq1ElwB2JcuC+lcOLRdGrRPi69x8vNnb9ZICp
G87R9rW0XgWXJRdAI6VgZqkYVhcTbDf0S+6ilAQH6x8fj0o608kbLBH1i6BBa3cBBrI9k99/hltt
HfCiSJQn7W9fa7qviNFtF/7xrTTdsVbpHj72Yvu8SU7DBXByPa6/1SwsXbbC+RqbfXzDD1nPvm/q
iHd+FW7i2jfdrYhDidd/xGP+jDBVRyzTH4IxjdSgNOmGct92DRw6dS5XaYbAkm09JosrfpEc4Ikr
hoTRsphgeNQ1YGUoe4JhI8RRCWeRcSWS2gxk6Ncn9wXpMFNx6saR7PjrfmsId4IKHWr24BS9qXcl
YwCn8j8icGIVo6mk9In46yB7LhBFBmQLtx4uL75PdeleMkRiU4UbzlJkl0XDzWXW3fKmGRCEBQ7i
5AU8MrT8HgTKQSOYn9+ne5XRPd8WqQ1HophHMKxTJHNTwzGHqRDMWzi84wjLwUix0EM3+L4yN2ou
AcWQQtnsE3mjP+UGmGg7UqpdxAJIU4uYSouD6EUHolCUKwLMuYPZ/QIVkdCmJUUAkzJ2aEyZjLH7
nhSZF8+YhmR5DDx9awhPjpgseWBYnS6w9VJLBAtDaWwsDJM3Z4cBqpb31gnoxr09DCwsAOxdpIZS
jvC/ghC7HIejxO55zrcrkW/MFKrg8ONVTlV9m+oWocHCAhoWbIgeOLdzDNMJZav9kGguVAtMwxwS
YBTMcUwKfbYWvil/rpHQA6PnlsE4yogaR55UZ+sSg5nk2thyarl8Er9mZU9cAiMapH1vpvLg5FMf
B9UwUcauadDAJ/8QA0rm8nTSzE7RQwmf03fhTidnt3CmsyIEh9fUamYYojtHFxzNvhpMv7CLstsm
HEchbihdeiqvp4uqXEenXspikrXoO1gMqOeU5AZOv7M2TI/lWoCmEfa2/Tev+2RpepjzpOEC5u0w
iHz3WAvt6n9lEvqiLvW7tQozjGEiOrXLCdYOZzwM19lv/M+8b+16UKCvqQnd6hMwiC1eBABMTxH6
iyhL4MJw0PeAVrfXXcdzjLGjtKLpvak4y1ijJubNAd80EpQMs/i64bKuHAOP0sLbgJ6TJamp0fML
9aCIM0LMa/Htd9iZEXgAQc5vs2OH1nN2U9jH9OvFlMrRnSWnexdECN3xE/NATv+T6Adtlfc8lU/t
l9pLHAwJ4e/Zr4/6GgpwlaEWRWtswqsNxP/Qniu7QWoAjjQ2UmpYs0WiTenI7ID2RisOqP5EARlf
eQN4vIUiZAKkHcg3ALXo7DF77UFdU0tJ2/EAaKRNeYaBy9ib/PzVCGi9a0mxJpW58p3EFKsxZcUS
9UskKcnXvwRKeSlc8DZvGmN+EqxFHf8nX2XoMKGSZjzNl8ipeIx+3gIvMICdYNWP5Xcm63ZGq7Zo
fCHB4nh++yZ2Wghu5C50vWQNUDmeVCXk/OxDNLcgaum/kO7WfyFf06D4POVIrS2tvPbgwB2f46BU
KQIBhhR3/YwKyArjw+s6a23wpbhfu4KYQix9fXIwSrrKsuKkaEc2eX6N58FbYkq8Js4YcANjJJAy
lKfecd0oZoI8G4/79VqgUKGG02kC50Cra9SsLhhf8LeTbiBDhPYuG8Lgzhi5u+gpwMyTxFXGUfqq
/F+W2D3mAKZ9dorYs1pSZWqIoNIGqh6dUgqR8cAzUo4R8xcemQdDUmdDx0VfCJJ2VXwhlPPbRdFq
CBxjOYXOT8XXejNdf7a9t2TiMh7DFN8bSQzGPtsnLN9yH2vsc4p+A1m5rLWRoorNc10bGDbuiZGR
uMee6uP3+d+urQry4y1zvqGaB0lxTI8MGz/un+8ykLWc6InWzvJYTYklQO+gbhcFXaSz7Uoj3hYo
e9y/bIhHKzh3y8i3icZ/lZ/CHNeaEd4mOPxfvx26mO75AnXkAwsgxICO5D5xo2y0+ZRV1+bBoEx+
hESp4qsrBYGnO8r4KqtJvfn2qjBGhrz9vGNcOZ7DVEDFTIfObiXNAmXgFp1+HZcghlNXwa5/FZTZ
E72g4pcU7RAaY+qWA7wKLz5ohzLjVhygC6OUXfKzHjqbUnxAsiC3DqzmUvhk5NC/TAXt9+lQUZXZ
SSmHFYyzpErYsNTGzUeOF1ksO3jj/iRXC0DTEGrFWKenli0sE6EPkoZ1gyMBkXeLe8AS/DSKc/D5
h53GotcqddECqCNnPzc0LdJ4FGrioh0Nwx5QqImcmer9Dl+dXxpYYLkR+vTXacsEH7m759df6YRY
IMoFvwwecOnafeSDX/7oEQi+FfVihn055N9TWTBCD+r73WjAGq02nCqQ4J0EeZGGEH4tXTzsU/Tp
Bz5ou1F6Jd3kZ8jMvxMg27Cv+LjDnMaeDYuwM7nb9Dpd0+vKXpeIYCGpZeLVmATpJHswaF+TfzKr
Io5/LLsS/W9tcPj+eRH/6WtpDOHM9jpdq9/hyEOOI+f3FZ6JbOSR2purHLZrxvvmewJgWmPK1RHL
tEwv90vES6qGyxQl00jliSgr4mxo2L0Rns4B5h4J5dLISX5npZx8qTMPBpnPgbLtC8T+xvNRZ86X
Zg/8pgruVJPHk+36g5L8/0CsT97qMeAZhHvkg0dt9DdliNlxBSEP4SiOj1Ng1HDPnzjC/fnn563P
uGbNg0Ar/jX/jqb24AyicnlDZ1PXfXlzX9Ikjve36VfkPApsOrF4dHd6pKkJsaeHhxMZ47c7O3s9
2T3A1SH4PooO+tiiitIWryACp61XFQ4E+pdHGdEXq8bFsN1H8XfawTyBAgJsAvB2YjKwDs1KtBvq
xGAOIWDXZBbeCOcdhMi+eELTf7wqDfS1CiZjhbAxm7Pg6scm4tmKLi7cYrXM8kEWESBPQLLGnp42
O4YD3oKvwJpRORV64lKIp+R5wd80baJblO7J407UuDY6ceBFWahD98ZeNxGkQZi4CP6jTRi+odjD
8dKG6qsRbo3zUtGWFnff3taTlgKGGIgRK33JyoxVJaaQ+1O62vQKEvXi3cDni7Huz4/575qw81rm
U4gy0Xu0K6anxKx+AAE8OO3VAyKbFyyH657u9xe39dvOpG6tbgdyIxrXdJIf1svlbVK4KTLq1M0+
i6mZAnBjXixR3Qnq28jxz2jFqQ7UhUTSE8JfxQLHvbyFlfolt6V/S41coqRUyDVRR96D+JGrwiXC
guw/oUrNz8MLjwJXX+lRI/gmanB/g9GC1nSHcxn3ABNunmoTIGfN9pq/mprF2kXUsDFO55M17RFm
4Wg/l5ylWh6ur5xdqDQKW/c2T3Rs93iVdf4hTBoc+S2II0yXlagfHt4Mw9AtvD2bJVmt8JEDHr45
mbH2OezspWlKELZtdGWPiip1klOlGv47GDoYOoyK5zIqwRWhtdb1DiQ6EWbFz1Vj3bYZNvBCnZc+
hLQtBrNhaxQHtIB9PPEDgTJLPS6i7n+79CQ/j0culXea6PZ/dWoZPx1mnO72MgpvR+8HfUCiixF7
QeCms9+DdiaUt8Ew9Tf7wdXOrTdJudKJJ7Zi5F2vacj3984dfPgAfxOGqw/c8TeQMaXkAmg7NtF3
CRQFZ6TR92HYD/ZbeYSoBXpLX+CRLKkPxPVCeFye2zdxX2E49yrh4fR7PnTkRHJZf5BZsOTtGSc0
Z1eIvckHC6Nwf/9+sYJimeMVq5D7ljbEH91JPkgN/KyP60dK8UQR2WZtD0jKnek5eTShYmhbbKJe
6a4gMWTpRTr2qViNMeUir/J7MB69TZgo4+USgr5oG2Xgj5XiPkDuduSKGfLToQvqm8BBER0kNxCv
6n8aDdfbsJMlt19DuTYFXXfF8JB3XRFGXwA/jInw6XVx3JZUTSrDINnzct4NmAAcwjaejQwaOGQH
ucXYy3QmiwPxwtQRwMev3055FbbHvgUuwYFSIVW8D+MJwmLr4eTd09VW1ShzzMLNi8hOsZR396JK
AMrGuVwCdEMzJzhdCydb7rsb8vxZC9QibZ9NGVj0G0FyaYrEFxWEC0OLwVuHdFfjywiUzFKxfO8I
6lepeYM8wNqVomEw4nC8plyR8gp62ViL8JOjmlWc5uDNa/9Qx7ONFcdzzvlV1WlfIk69b0LwgH07
HbGpd0Lo7kLDW2LBI65iZYpb19hMs4rht1894rx/YtQmAOm2HD0aXJOLPbwP3qn4JaD+T4d3Kbcu
+jqg1PLPacjp8FuL64pj9qmr5knCBsNluJ6vr987er+BIvB26LPyUt07G8JCpJsKKRbrcKUZ2fpZ
UPaMjP84axfqJFqeqbEb7Aw97Rn3jmX9RyH21rB1IvQ9Pdy/iK0q2hSFdo10t/HSIrbEK41YW+cd
uF9DB666Oza0z00ZoJCxhkhixYfW4tSur1XXa7Zw0aoMX+f46aeWMbiDWjhLf7Z0ez0WT1xLUQNL
1ceQNj5OZVz9vhoEWFl5x5nUAlxwN2yMC09x30uyCZqfU4pJyIYMJShJrpbTlwQSeAIYXP/3EdRc
pbLvanxY8d6yMGrpOAJwlACZCK6/F+9Hhgbd5UgeGEOnqmCLXPwaTbl9H4qdE+ThT5n+dwhZaSc6
jKJg40TGyrrwdkkGR7PgtIB8jAPtXC8y5jowgsdrI53iuN4P7/vlmSIGg4jAIKDpPnyLMaLSvUcu
ZXmsUXW/7wRr+9Io3iMYjEFR6djMGqvM3I0JoqVtPr033k2Un9MiUFVe8LbOHc8DujwPPdrBxM3O
I8gCl04uyweUuwvb40kOCRcxuvnOqPEF9Au1fpBbt+Rxe8paySyqLcFXh1mN84l6kepEL0aQ0Zun
JWWj5NWVKAZrWMqIPSTZ1FAidRA1Cdn3EueTBYyRjmrrdq+aGF9h7XkciF3YFk/Yi4IlLE6NpO8U
7oj4MKd5serRb1P0xWOU20NGfqvIRW3+BJeB+jweSBN1/cB8lCsjBPQ7XZyd8eZxrMWnPEEaIEZQ
jqwcKsjtZpyC4MiE32QN0eCNyI+S+uRTcfqRFwHcpaPKuZeZ+hlTIiR3TVdKbCMowZ+Oafdn0fNA
sBfXo7jinJJdP7syv4v5na5IxJAM48wIy3KtLOYLQnOOhLQljgHqxfwbHQ8QC9Hdkvpz7UgVvYCz
8IIuim+8q0AnWurOnz2RxmYfF39nsL6+tioR/pltg4vu4OcuyXEidGFomNh+71LtnKqVyOg/KqBM
rqqkz1lp1eAXz5uOg2eYlXsiRMGRd77TpBRPIsFUqgagDBCsz2Ls3U08W2V8SZ1oHrBwQcL1EMLu
mZHhapuSWq/LIyjHxxf6Fb2rs4YfsbiLwrr4A/mXqBiJCntKQlkYK2QnP4P7NPeXHk5THBkFydgp
kP6FJQ5yvwr/HJEG+iSelIe4E51G/fh14XD/oZoM/yGg/Nz/lyMlotiTUTHuoQbQ6cVeayV82ekT
XYyNu/nubQoO8oxJzflNaC0dhqR7luCOXcONQBi36mDTfwOZVKet/7QdUTNBNg+CCEqVvVyjoFBy
Hh53qTH/iE3eOnSkCCO8oYaAvYXjth4sIYDFD7SO26vVaeFM/f5QBtgaB+xTEUMEum5TpdZ+Cn+7
SR3VJQO6JJ0wwjXzK6JL0RopB8OeAa9Fr4XVGjienIUyrnDzkgUcZdj0GIfWaL/wc5lJY2ogvo4S
Ayq2LhNsaGOYrZ5ihzgrlsiM+5JuI+xNYEsv4ON8t/KOS3JKKX36Sw368K54+0wXAXBXHkPWq61m
gpddcmLd6e3y2KX8M3I1KRwprGUoUAam79Sj1VhMVvy/tQijo2e81EJd3+d64bMaXA2pfQkT+K87
B0erUzmIcwoRwMDtuJW9/RpI03nIfO/CQBZ6IqAz81rM7KQuhjclImPo3WNglLw+27REw2Dlu07U
cMHtIwBDzXAI03Xi4Mwij1owiErHSbIHr5vf3CtglmEGbwjuWp2ItD8MTDKYKLCVH2ZGFLKJlWbS
0gike1VX7Wj0Ay1lo5jzlxWLiYZMbc9h28F3UWN+4aV7xwGL7mTOp3JA1IP1WwqR4zAH4Txk5nEN
rtppVsVXuEAjp5zrxK/jXlcmamSyYXCV/UREBboqjX4maxVIEWA/kN+JR6AIJyKK8AauF3uGVT6q
+zCHldC1Xc3YO3yaP7Hqf4Af8Gnv6y0eiMbzGjJ7mSdmgB/pQ5zMfFaWP69uMO3GYZkRQtV+lGpr
1ErXVN/j+yu5DMdBGApUUYeSnmjniyzt7sw3RNz0m60d+vvDWupFtDD+K1M7katLCPVVzeJKP/g/
b5nYznja2HnhFqwyAheT1Awq/ned6rpuOk2aglGI0QzIvICs40UUHTYrCKk2lhjsVEc5zk6mD54n
kRiwzrof9Z/pzNBRyTM5V9Lz6gQSh7U2pSFFJmI1RO7ck96q+wdcQxVw7zpPOMiCYgEDHennsTGJ
RlT+0LBZ+9KnPWW411NvLlMWWWrZF3/hUZFwMdFPe8tUelwakf9vcUFBzHrtEdf4UK77xMKVKFlm
aIeO/dCRhvOKDoolqiQLTLJpNy8rwGXmTGHmivLlDJWCB8URI5bhP7Du8tC0zP0dXDxWr7gQyvQ9
/+EB+IbDO/z/skyNN9W9gl16kN9PjiH0F1gIe15sJdzIPZny30VOMP+vGTCZ46AtKmkxXVtllLDv
rKiZ9iymROG1d6D1gI544P655RWwSzh0jcmyfdqSOPiS+RaXB5m1VvQd26/NRtvDUwbrhCi4uTs9
VgeDgrpHkCA6F/cXXP2hhJpyqgo2L9rMVGParyelxaTvXro7mEa4HJKRVPrT3bg5g/qqosLWA/pO
BVOGXcKpsGQAfdzKdCRd+ZlsMoyg44WkLG/Y5lyYKIi821ORRO5Ldj4xBkJAc4tndp7kBcdIR/AN
RAgUcDlLfjKcCazvBei61f2Mw4DGuwbajo931R45OqD5GHfzTRLs1QcfFy8vROLIDQyZg2R3WNdk
fnCTSlmsWP6TUXjRv2hwUbWQz/eD2l3kKL/gLVelW9fvk57sZOUPuGcRrkvF4yq3Wn+nQsM8MLeQ
3v2fA/iVw5AfXhhiGq5BH2EF9uiiaWmJ+bXcOE1+0ODSQZuos/4skshUUIn1tDsk6tFEdh0YcwK9
nvUJDwuurQgV22SRcI0qPv3l2ZpcajEE98YwconA/ETFFscMx5JnjOrl13u8nxFFRvjJ6HyrRxPm
IwLG80q/FLMVxj46nHdsNY6XDaJb0kuDtWpXMUFKvPBdiDKRjNUbP2uLfQ4B7tMxc+IjIJCNyRYp
1WOrTuA+yqmO1xGPRYwM8EqOxXKpnuffGBLpd5sgGiX1R38ZHbF7oWjxuudBbirFMxYAlRUfOkrQ
3YfEykhBiBGTKTm0s/xMONAKeQEQLZCHqgUbOX0JrnwjbryzLb+sMozfOKrG1pLKItaw/u0U/g1m
YN7yei8ajYK+rkyo+o+I6MkjYBCXQH7h6jok+uS+UhaFF5nhjnMye7pyCR380PIMX04GPX/2ICwK
uTO6QdMR0Wh0i6wHm95nW9Y3n4dcmnql2gxXRaSF67s42Yg/IKKEe5v2IbraV7VIPUTwhLFlDIGs
Yty+R2eq2qqTYz+9ZSgScqz/w4hY+epwjnwj1e/zaV4Zct3Tphi3wDVk2A2RSp/f4FBilVdQGxuR
GmBI3c5+Sfzd5dZxDsA7h2QnftrrKTJiIN6s4OyTicwpnnx+aar6Nw01DdVDKmpXsa2p+/H2phbK
+QOQyOw9B4HsmpPVTHW6aoLi1dF5wtwxThTuEx0QukAF++1b8WcMQXBtLNc5Ao5RtSktyH+3trJy
ZUiGRp49AjjZAIbB+Sh2D5SGBM9VD32CLJXeKKtmpei0vanWSJI/b3lNB1hhjYVqxkAGBNvKkbiL
4UMqzeFu3565UfGrTVN49GXW/WnB6yoDiW7SsBnXGbwV1S6mez1R5juEZjEMjwQtTBEVkb5x0fLX
VpdtgZYleFMpbwBa6Z1yltDQfXszPe9rmj140UBsJOmawway0Wz09jCKhwzx0v9lgs/YUpgezbvn
FI30fwZwnVtUnR8umU+JjUEiQV7vxB0i9VT4F+7IUIpD0C0FvaMvEZLaso/GgfVMfqO5s/GZk+u5
NYvlVGoYX9kIuiMMuP9+oRouWfxC2nYEGI2TNV/3R1dOaiIEsPrYM+ZRd9dISyAszu35+Zpw+K9r
Q2HQsI/toXfkL3wqqlZfnzUxzSetecGyxzB2hOT7svaBKSZWQq96lP26jjnKVovHIcoRLB1AHVwQ
Y3y4ssvBeuNrYZEbzfCYspU0sK2X8Iz9TQIafizSZwDUbuNEIdAjx+T6/pIHqwoqeL5boYtxrED9
PAQThxDOjMLYDm/fWurhoqlKbz1wxDP92IJsvlRFfAH4oc2z8LnAeZp7zZnXAdZ8YdshWDH7EoIC
gLY5NOpj/wBNcUpqrGv9NTMo8Pc/FzuSYZu96xjn3ppR0axQageVJwQI0olo/r+3VaQ2ha9WUTso
XNV7lpa5JAoB/DE5xDvI4Z356MvHCo2sFGJwqv52GK+Qodz5mCaC/H6NStVEefWGGV8uHyTvApa7
tIBf6AY7yhtYotBxQQ3Mza3kyHDrsZ5IrgYBEiZtjxBMCJgEUuzbnX5lYKK1v4lwwB9GhVEnotOF
UjSimVHdoMpNVJGda7mOfsruf3loa1/jBa1vPVxaG9vRZCnH1cSdFECzdZ9nh//QVsLxHhWGbeXX
Q35RKd/bj0Q1ufeusrUc6JaVMY4wgi5JH8+YptSYdao0PMuOnbNHiCiG0wsGjnCaiGiwJRUynf+t
Ja1sLgbuiVvjRLiifWxlTz3k9HZuaxKHQoRepWuAkRMs2yFIsCaSAuzRsrRS8Afjeat7zAgiIAIB
oJJWrro2uuA6wRVL7b94X3VMaCfuT9VmAqIPtwj20EchUYoLzCt0oGGRXiXeekUBonsAXgpxDpEX
VJyvdf3/u9UdMcRGkGbb4UITZZ99UjUpT/nRldN916IPM5MJ5JHcwOM8Uf7vDlPB5Ll5ZwdkjXWD
xOznVe5o17Z27vEbfYO1pHcYHywUKZ4+ReLEKI5uk4SVlM+L2QCZ0ieDmw2h3XEwTxbQBBe0iCJK
kLAEz9nY1FVl76vOCr/qYq4gdXCKf1Dwk1IaUvJnjY1VAfEHtTQFknaCQdFLXuHfeF+xAUVZcTRN
fo5Y8lWkzyzaxGFlVr8/GfrVn5g3YmRd+VKhyzRXML5iCWzAzxrK77SiFL/N8j4z79aqJgTg2ePH
/FKk9rzdgqTEJLDFRkuRi9xdyoYS3bnD/8Lx703Zx97iyo2PXYSWOmC/Wz2fMOir7m9f4a//HuJG
unGNPazEilfcKghQCHYOX+MHJD8PlAPv0wuX151vYsgbcF/5ZI9a98/zsiiNSWYsT1xdrRhbDTB7
URWXF/GFqtUo9yXkfQ1eHvS6+0NFMXfNWA2qBmXJK4Yksdq/8wWIBHl6fMGP2ItfMHjy+H8/7uXw
6FbksW5a5C97dPUTqBPfwR1v5I7FxhiThNE1VxosQSBtX3OyAryoID49t5ybxoqaItNMD8J27aYb
ZPG4RnxWVGF6wxJ/zNHKCY0jA8A3q0HoEmxgQuaaKYMJZHi4cF2fjv0sqft7C2dWL3zVyF0RyEyh
WFnObtnGl0HFHIr8dpfWlazi57IrEL37WwqIqPIk4tU95+ikkkwkbl8IgIh+BX72p5ky/OUoz/oU
wGSGeUkFur+lUitbzbKsHWzP2Aw2jdpgQ46GykWeYRiSzls0x2D+F+GHs6svIMndMxx+AGQUxtTb
MwHCXWkpHzBVZhN6uOcBpx3WZUP8CiMQZTDy/HLUiOaVDtMRYmpdOQY0wWzwhWzbXGNrSoEBHDlF
FgSbVs1jB0PrZNmpMb9Wm+/zkIKIYAkCK67pIgga2XPMf8WrGOR2bEB3hj8/QA4kCjJ2HYsgJhgY
qcPSCwfr2WmUJciUXVA0Z7WzVl29ff40S7Xx1PRsv9BgrXBaoNGlb6L9Ylc8FdC8VjOLYQEJBcWv
4d7YV4uXiavykzPbJSeVA1XZi6KacTcwaN7m9D5Vrie/kvGyrR42LVhAzoQbQGTXtyq97LTzyeJQ
3f8UvGCxGuWwy/U2elhHXRcgfbhuQF5RfVtLeCBOcNxy6FqK5hrxAV4vdoFY/XXrDz1mpS0HMngD
lCAS4vB1BWH003xLtKbZIs9TDAuZPy5cU7KYLuc8vsnFDE/EEiXQUQ3o/ZTt5DFZDkHwP3q9dpPs
hbs3IOJCA+t0BFAB+5hlmVr1E4ZIC4+r64gQwR+LLhbN8YJmlYZWXyZgHsQYLy9fneUPRYMHspFA
jbnyv9KSyd65jE1KlMUIokQnEUoUkQYbUR/5mjvHTXTrRhUy2QzI4PZ4pEaaU4U2SNKHvjLCBMBW
rAHWAcjrm/RySBuS3No9d495eotojP7OgVu5u2jHmwhMCpA9T748oOfJ30W4nv8/ulNVqts22jRl
gtS49sdi4QEvVH9s7u2i+GrB6ffBf7h5ZsfyCh1arfDho8wR0fENQjrQyhPuKcRcSDegSDU+LYGF
y6E6yRKnaWYF8CRjV0mPy0oz6GqrL5fmqLu2yzBNi1/X0LFvHxmF7JT2E34+R3l2yAqqQxoC7LX/
2SM3ihyCwYn25vpldn6j8r/rnvoLl+Nf/40p3MLlj2NaGZo/fMLfSrpLmPRzRvhlGKAk02wnFrl6
U/D+Cx+71O5Qj0Np2bKvM57QRyfZhSc5wLccdqziwiYZnHSLtkehhal5xW45ljkDAbvdhANzEgSc
Ac0RyDWekpjIofzO2MH7BwqHq+K/ovZ4E7S9+oeqcoA/XnV3DbF9IIlbJEpA43QcSKKTMpCgzFLl
CMMLiZmKydvurrbJtcv5CAFbobDoR3Bs3CCrymiycR5ImOU9eaYLwR/YjDWfG5BatEK+khPnc6bj
cEU8JB6qfLY77DfQfotPHo9YraSEpJs892WIBChNtw86y3pemEJqAVCXnErhslaP7wDv3VDRhsPX
ToeKBbTEhpVyycfVY1PKJqKSuGKVlpl9i64keq5yFgvYZkBBF6kNLUZGTwgJExtngxpUux0osBG9
OMUNGXSXy9uFSGmnPjuP2gn9ffsaHDK0PsCeKTDdfa08sedyRN7Kfp8aPYfBf4ySws2RuGekLck6
DFuFHR6j9dInG/okcgPqc6/OD3ndQ9ZSl2ymfPdmcbuQQ4PLkKl4ZZ684AjX9yhFMp2oLPP3T2vY
ILSA1iBoJ3mjHZ3zqs75/iPQV0pLJcwsH80OJIc9WotIMKftIhQBnWgdWZDIhHrm26nKopS+pHs2
GSEmYMT6Mwxmii6v1etSyJairl4JDXQ2y/HjLKiiXb6Q9prRl+cV6P01Ku5nJeMIOKr74OhzkBhi
Bcl5C0mSgFXLZbQ31Ow2F9HOxWZPQc02s9aanLPllAd7Ye/qB+ehTzVNqfp4M29QOuoWccUBFqIQ
ErZDmlqVD7UNUxEAYFrMUJjEAaHCSLk4mWpwD/6UXmIKCJC3A9aGpyHkr7WUZFqXLzfkF9wN/uT+
8FRnWN7BMrO1Y6hzImBp1i+iMbLnUVEEQFfhPqn5vE97jMWN0EnSNzsec0l96f9Y91tS5Aka51Ay
oVaLWIkgW/qlNGCdRrHiiGuAVeyYoXJOHhMANObihugv+ItkMP43MkKT66yTWMKactoFVAGwhydx
NNRXBNX9OP4xubNA13CuQD3iusvmBQQtNeA88Vg82AoV8yFelimHjE0lLfXh+8gXT/3KpiMo9Ab/
xueOw4QL6W+iP7pdp2OYbGfxYqmpvJphqW9XL7AJKKSsCh+dS7ZuNvIIWu+Bn4PcdF20KqZEnPkc
Ln4/yzAOGt7kGu8XMn6x9QI6m2BEFYWWagVnxFfwtK8RHxL3BFtQonMIMcxGSPzUtkq075yiDJdZ
fbUjSJGfA8YVjOUxnm7f474uHRjdiWMni+akNGve6tK00oMyEznw+8/IrG1n6yBxWdYjPhu8DIWS
3dCixrRYNDjT6NjTIxPbssVrofBlbrMy5ER9/Sz0VrVwm20H4mfQeSMsbdE8OLwFrgVgc/RcYCSs
t1cWF46phObcthzv1gSVFoqy6iEowxnbZCtws2cWcVVOZD0AxMimZoVwAllqdMvcZxDFePexD0x5
z8kCI/jdM3dvVcPe43gpuAGnaN7qdLYlBxoDMCZdvylsm3oGjAabv8Y6g0CU9HPDpJH7fAlEowUk
RHQTZ6ezfC+dEEY+XJ3ADB38yx7OQltmSSnASlzf9iuHipus5nwVoM+HB+p8pnTYTDF18gn+NpNZ
MAjfU3oyK2/4FA8F/9dI75UvLyRP3sYqHrky7MAQd5QcO4C9BF1hrNunyp3vBdz4+EjUunXRMhE8
Q8jJYqIexQPovX+xGLKYoqOEE0bxFFwclUHrJr1EgdU79IyDYW3Y122vWNRTlFCghW2ZS29gkMt2
joow+ZzXyhpfpQtkg60UY/1KTGeh4tEFGtr9P8cgP5mA9fOAW7i2bGR7rtVBKoG3ixYFnCfQ69+t
aE/KexslKRmwpkhGsniRdNnJ+nWWEzZHglZi8kUEwGqLs1d6vJSj42bZs6oCdsB/IzY5wkUExgKg
YOaV+meHKI1D3A3cnFdOA370yniSk2ccNftJal6G+OZtUS28Q6ESaJHqVVIieeVnbiTdVwwYlBQ6
EvC266XnljgP4kRZrG5QSk8OoU6MdaOFeNHVMC+NuFwBcjBn4QOG8b1Qn7uE0Ah1boGyf72xn7bP
wx0o/PR1+8sMAOvd2hHbTy/TIqAAiXoF5r5bICi2o2nMm3TmreGDV3yIYZ/HYoO+GOzx7ml23GlB
7RBEOyoevd4OQpLq4yfPKXi5Ny6dHWyGR6CUN6dHuqTLHHLzXFoUYhoEK/YkBiMrYjIbr0qTApQd
i0T0/fy20zxEu4pL1DiCX6QL0sPUaNAGF6+IA25tfEiDhq4I2Pn5CKm4uzRVYD7GKvL+1Q+060V8
qILjHBPnfQeKFcjTq1xegCqyHvWE+Yi/yeWXj90UTyqnz8jGCFeAPrs3Mm/NiIY0C+N5z0ZmIoHl
ojwahZA09dgwvtu9Aeq+mOLC4E4eK8ToZRG6/fpWOAZWauC+FGH5Su2P+WAEAsc+Vs5Ohy9d8thl
8LrIfq8DH1p0qpxIub77CyNC0MCRntOEQWC8b9u3VwsjlpjzyEWGkEXFAvoX/y2jlRfbD8/3vLP2
ByYc1x3VSt8fjW6XGsLOQjoDoIcEAYxiucmQX0/7Vh3Py9/N9yttVlBSSNGyM2rtll+TbALaL4jK
dqot9MNKWbIMf94DOGLzI8kOjxqsVWl/90KBnEHEDghjqIYOkK//CBhamezkr4qwihAuRI8ZxEjZ
yxbhKP4+bfMppZVm1EqyJ6iJFYOHt60pwNGAVAcOjd0Ab2AkAWTxkDWDWk3Ij20hOPhTHRFjZi0c
9sQiha2Zl1NlmULYbwTmOcgGOpG6MfNPj7nQXMon8SNi8pvQWZdZwdct7A0vcPTf6kmbwrO+afJs
vw2nZJCDf1RW/TemCXVMlpY50qjDUe/xCeL2LIig4ozTme1kP8fncl294wh8xNB7N6ChN0Ect/p+
qaBy3LBwC5tY4NB8FwEBEPv9cQwgnusCeaNaIfdKI2aZA/NaSx78O65Px5GTaJd4uEceIh95JFJp
mmG3XH+O88JxOQb3AaH00oEaHgpEcTLpdVIDrqhL0lhnw9+sRVGFek847LicxOuYoGkSO7XB5zZV
C0tn2Vv4JGTPEQ190wmx7RtDMMn1OJAn1dEV1HrHVqUud01t1ZrZPeYEFlL+RyDhZGYK3GyRnhid
yAaGY+eKYNSzlnoOJMyQoujk9jTj3g2xSledoFZ7R9YbsYVe3eL1d4WqWjg+eSL/sOMJcIX056Ko
N7AXjw4rDnP7ZA5+NL8WYfbYVVIR1jDxAioEniYePgb8da+hP8weW/ipZWRnvrB/dPhVhMN8pMYu
IvKdLln6NdaEfuicmqA1b1TlTWHqAMlgcN8shVpG9aUxabV9+eOWD0YTS4JqGVSc6P9/2Plsc0yp
915Egy8OOoz/ovz0GWkoUsvo8YpSKF92fO4oPVs0z/WX6entkwfazSGgFy/P5aCbdx6fqsjTzfJr
kFQtEFwuq+d2kGnw0EPhnT726SOM4pWU1ghfIMqoDbbV1bA7qX0cb9H4EeoEtkPqpP8k+UO8uc50
KjzJXX8YCtc6FRp8MqiF0DPXFlSeAPFm4UkbhMfzrgL/j1eWMdRWq8B1QepbK1wgwpjk+RqgVwwj
Hk1BrzDqAXWMOuJOydpcUOHy5B0SOcz0dbwSeUUpJUMmZKq+1W5WHIuG/bMsA9RpQf9wCmlZxu90
0eKbe8qfJc0KkPEgWJl30Xdng1+LChPnPlIjLAmqxQx5ZIGJWIiQIUsdaDU1B19SP8eCIoAZOgQg
47YqpdUJVRxCoYoiMNU5deZvi6v7AxfAjuCqmZFGfx0/gyk0RZfxq2a+woaraUMccq+kCpZxY2pv
j9oanr6mVauu3sVV/hL1X+LAJ0sg69o7G4FCTZu8mf1aRYYfFF2iokf9z2H23alXAx4rYFqT4rEj
aRB47OFp1DS9z6cXK4D2ngkM7sdZ+u+KuH4mflzKNg+mGDrTm+H5N7JAQ5VtT7wLMA5yhWuI8toX
1NrbDBQzlc2/Iy1yYp6cOMKrarjNN3u2CuIjnoBRAC/63rk3SSd79unFKMGkD9FYPcYnrbJrwetk
3hsDaphEWXSanoLEUgFm4GQ4G9f9TDCank15/CIDzNsekH3zPNlGz3TvEoY951mErx+shV76FyWz
vhJ4OIvhoqJ3svC/aPLlUvj2jAU1CqhR0yMMw4N32PUrYD8RfuYz4lUBfC1VsBBDMppOyviCblo4
wV0zPUR9P6do/8/2zmNcOmjwzwCLRGZpCf4fIeGgJ7scl8AEh/t3BO0OfIt+xqQiv8nfrxDPjZ+a
kvppcbNrz+eRTwdLXTIyRdC8DAyEfpMrsDd2lqubt/HJfJ2WsSVgv+6ZJ2Z6HXmRgPdxqt6zLaCH
OidBOZrlTEL624M3Anug+gpkdH8E2XHdgyYTDuuRIvsbBIAwL3t6VTtcumvQ3adbG//qMTXQR+lD
wbG9NmPqsg0AdSIHdJUaWnfqfNgQn+xsx+ExR2OP/rzSDF3OdBw1tKfZAF1WzNmBBz0Q0G5HTux1
OggvNiDb3QQMwmyQTKjtNs4uP0xoE4j8/XUTD+QONPRK3sx2j4N8GpjADrq/VrjY3yp3NfxDYUNy
UHTt/jO3YUEf2jJNeh4jiCaYDCXj+S2VDssBkyNGBmnbfS90q2+ApzuYV9UpKJE+dxMTUvKQXk10
aZHshZlx8UwhcUnc5Pq1/c19VSuDeL6/nF/fPyJLQn6UxWvFGj3OVcA+luNUBo/L0iNOEr7WTnsd
ZMUsA2ZSN2csEsBNvXiN0rlZYzSgv27UrQDLUNsqcNLyFGqilnJcHwOotv60OxZZiFZvoh7Iy2cm
JMfiHo4yT7xmaagnMMQvdGM5ZG+j794iQrFvV+KKH7RW9tDOnOOGgQumRpKFSOO/H7kPTgzsa/aU
J3mPamScOnq7sqiMVOZzgGQQsGcEnghYMUUxw+nD0yGMQ02FVjCrzcLpEj0MD1eBL1mNu6d1rb/V
0WSn8vQlN10lyCKZxac0UD10CcHJlmrs2SYhRgR4DHUgHWvbj22OL2/FxFOu2xW70id+GaAA64wm
2nqdhycJXv/BGhNee08tyJD5KDa/L1I59YgS+NB0Zkmi2i950xsw/FEXAaQiPf020bLI0g6R/pP/
QyEQZEdc5GtMuxN/qZPvn+XfiqRSvPJTqJUN3LUBV+mpuuPqKnLW7k4iKIsYhEwHzQk6BZRIMCJT
4tvNZme6cgBpBI4BMwZFBmRu3seTab8hUEhEmfZ4co6DS65JruvDk2oIQnohir/Gscztu5VK9psY
7CUr+tcERk4sWxSKm9xgpQI3fyj1RNPezepEa4JifQpYbmOPAOROnqEto6tw9FdTah0wlkzYN8Jv
6svANzcEHuVEBv2972DJYUdBeCRV5Evp6p0/AeUb4yH3aLhwDnp5EDZJQdKiUGvZ8gn9spHPERmi
01IwmofKRXEnAnbymhFVHKYTZTVVBWlTljmJaNcwvieRaU7XlGyHwwqimWRB3KpnlwSjQKn0aQPR
2oP1HqYYSqp2tlfOtiu26TyyP+sG+Wxk+ZKm9Of96f5gI9UqyXsaRdRzQ6ZJ/tSno5k6SGl8Prfs
4xbHaZNgYxoOdOppo6SczhY1jAzxbA1W6EG+9wW0Q73EwLCyLfR50jUaijPsLAVEMn2fEQOgCKXG
L5Jfp02ax6ArFgQjRMN5wKYiQToWLFMJfrmQMIu6y3MjqpX4ttKrLxRkAF+TYApah+YtY3tZ7nhZ
ANVIDvMz5xryCQsvAVuo0rwfarXcpVYfhxqI9nTgKFbf//LtyFmk2bmO4XDCC85bpZ2/pJ2rCzK6
9mpZfBx5+SWTm39ZSYzu46ojcdugYKX/YTN/dxpY5mC1+53hGVXewablcWLJZDKCS6R5cp/zXRQ9
QH5fSfD4APSAP33w7rcKTQatH63vLXFAR6SWQtZMJOiwyUoXOiViRpCzN9iXTGPnAf6J47JykbKJ
byFj82bQlNkrM5UiT2/DyFVp7RT2Hg6aBahzbhRtEs1/Tk2PTqbDlRuDOP+OjxO3i/dPfFI5d+Rj
7sMPUf/GLxhL+8owNLC2RXZxrik7qAPaTNH9DTZOvR8AMOZ2mrTk3q6oqoKN1ae8d1Yiws7yWRFW
KLWftmE0cWePyNW+f7leluEqH9xa9ksI5kFnKpRONZhuRoZS+AXiLHa92gvrJk68PgERrCuCPGU1
ESU6eeBDi08aGKHpJFrWCj8AvWViVYfdcoUwnGWSaEzzdjrStji9WyXA+CpHysXyt0dMp7pS2JRz
WTJfh5XhdqCs45kGDQng9raY29CZrTE4WJigECvwfJF2/9MkkzcPCo1xmwnHfhjixS3353ggmE1Q
gC3l0ArpF0lsZsTVD2xo4AAzJ4zjC1HoHcKAlhJm+ePUj+ZuYVA2d5NMM7MXnEdPJp2Y3ZxL2Nm5
QjHJ1r3caSs6uXY6787iCSmBSxXHqgTS24Zzyb1hEmmS77qMyF7kxqv/DO23mX+CjvCtOL1LmGYC
y3boebb9OGYKyjb2tSUQYnukEL7ANpPWBVH/OfZegP+o03BJhDl42u5tYFDUConvVo2H6/bB9zm2
hNGu4YMHTOBvKN14+1/5lrNV1Rc8XFkyqvTAwVgOITPU7K76PKEkAWoBGP6CvVdww2AvEQ1K0v0e
M2IR4CyBAfs3bHQXcQgDR7xmXP+FfK2gKWDcgfm9GJRs7uZERCK6M5lVDx+nZJT/3UoN/+8XF271
8VyGdrM8FgL2aIpSeAhxJ4gCRKicjjQWxiGnMQYWIPkSHHba4YFN6wFcucKgzKe1vw/1z/ooo6tj
7JrjbfpBexILFn0cldrog63f09XXZ4/2eeTCsHEMZn/Q9X2a2rvUeS4nlJNC8GKRWIHS9zf0zCGl
tf19EnM1Rg2FbA5eClUq4iamJzWviFDFgOwijx/RWd9vI0CL5Yu66TfeBkQwTci8Nlzrgl91+bd/
CpEQDLvJbPbZ8KTQRa0se1Nk4RSin9pNmuXEbVfvFAc46dkmUGtSlmOLVVcbtfmj+e/PrllN9pR+
bVxnI0RIjnNwL3nbPXFgT5Q6qlQGnA61UA/xlOXoXNIdH4TQDJCQaF+Cqe8Ly22hZFSh3bTxJzM+
OdG6IjNSH3/7Zl7H4/jynGeb+3H4cnls8ZN9i7bEClnORV9xTXEw5FkCZboVqNQhCHLvkCtTEJud
U/b39rE1C55dZN4Ak9xhD/eHrBpcHxixGToQUk4p30gSMdXangewLR2iebEK62zaS3HDttqxK9Xt
spVmyw7v8DcssdDY146AoYDfAMN6FAYEuND1Jw9NFiIdHJlTI0rnZrsnqg/u/Bhziz93OIcoDrVv
L9HJ6I/H+uOcoHZo6Pqmb/8iwGdQTAhV3zJIr0OGK+gEvRtYPNa0CbDicEOtujRnnkzSC95Gjd9N
9dyQ4JW1iBU0Xp48jYhnGlKFFrxmtK5CbjceUYl7tiEoGHQ9OZOCVVf2niiOBXsNP9YWBcBojbMI
m0IB/dz1vOozt73Qk4h4Ew7rwKAvGKLKU4UyfLyG6R7dpudbDU+GvKJAl8tJh3VWsCphXVZo2omS
DljNrlDmyeWDtnVf7iq92NR4xZ7WnNAKOMj0BdV3VBjmSW8KlupQY/weBA8cmfmiNkB3rCugHwwz
yXaCgNEWxG84gyf25HkzYbNtuv9JmhP703t2JzSo2zTr10+QlfkMy6WwY35QPxLnOMzeiavDQbyF
lc+RBz/Aqfk3achMgjWIj5X4smZegyD1q0UHm3cfli/5CviaE3jk+WkcdiBtqvzxn3TEugp+mRNn
I93RRf51ahD5ILI4QUDfsUxRHxSwLMTEgtf89csZmjn3EaIr0hHZ6+Fex+rFShYHyGypp/myOgXs
J9cRggFawEq/Nqa8TR4vaSCvSKN2n/zGL0rAwniV5byZ6Q/en/7K93BO1fSe//UQcB7VHfFUffRD
dpY9KDPLjrFEzJ6Vjm2QYvq96+6Vi0Td9/iQxAOpHen4InsqwLmjPUl6/rBnzI13dqDmBUn6vVh4
992PQC9+x6a//L2LZm3qalfxImabH7oJhNz2K6zfl831mHnJsAuzaubDteSc2OtEe6D5wYn1NBCh
0XIrrX5hAxPsT87noa6pMlcaCwXfEunDcRZfn9fyAz1rPwHWVXTzzrV9b9uoV8Sc7xX3vDq1yS3v
T2Hv4Mkjq0Hxnjcl7ORrnW7BGOBjWmumarqa07Bc/+Nkd65OgVvZjtRgI9W+O+uRJUW2j0ka9tA3
Xh3d1gyFeTd1RbsyEGCwDCjtpkInjOItt+s36mT395SsyCshqy6XJ9Sm+4XJj6TyLHVTeHhJR5T8
scoHs/h7ppXbVK+qR+bjsTsmSgc9PhHxjUNQd+Ok5aRPjTMkQ/x37iHBggqQd+UCZbXrckpQBKQe
a9OG/i5NFj9bb9ewiAI7FW0Wdg0JQezqact3IK2OBrp7q833CopgCDO6kUuOALneJdXL1NozqaTL
H6ynutliYekFZJ+tm64z6L69iDC14OkpcgqHy/FZQd5r6ODrCbfZ6l8fK7fjxgADb48+ssrJQNnn
zQFAdOSI9l0Pm8tBfLcKzBmFVK7Xua9F3sYNij/hYSjO3Xs1dPS+OARthKNSvx20iy2icTgiRxNH
RMjj0BXQWNuFPloaCBUaUli+m7jB7K5DtqdQSDurA+6Zkwn46XR9zRHGsQfWP5yTvoZIXwUgyO/G
SzI+yrjUWBBICVnDXsi+t4yAGs0+3/6RcSffKwTkzMpjiMMfT23S2ej7dO49/uq90m9iVSA0g8Bc
RXDbS86jlOQU3WWxcifK6gvtqCQtPPAecjczwSYH3scZx3/LCtcH5nLmbHaqKMhXgYrPy4odDLEb
65XmYh6WENj281HOe3RSM7Ne6oXvtPu5fUwXH+Y2jd2nrbRjCTzY7zDDk/1O+FDbz2lk2mSUrD40
ilN73RJ8wOd+u5h+DA98b27BthV2BR2CK7gcwzEgRT5jSN0Xj4eNHuQpt1GtOPBcIrE5MIXSU5Fb
DBgridBI3cwrLvLcLC8nE6yB9o1wIPisV7+p+Sb9G3C6kwCJhgPfwmZmGahBfKFfMlqme9eBtXBu
rgd/AXhVLLsxwjD5vZgrEhjVW7RD3spVTcZU8VKXKF4H96dEkXS/BZ3AxSh5mrslwA/xw3hil1wE
RRL09qZH0iZ+WZ9KDzVmYDrBPsHRcwxXesIV5AK0uAHT3RezygVghEZ+856jxOzAIPDHjG5htim6
XDcV/ZO4K+1Qo9CK8u45bsDyapMqwZEMHPmmtdv16FHiAuBokqZ7CUpoiwxrUDAef3PFqAem8LXt
mW9kTKnyU7mNWPtqwT2ej1/7akVhpMAt5XUhZAjC/RjtAPTSY+d+DbJi0CzeUgQq7bZif09Y/fPf
a5amKeaOFx8yLJh6U9T+ZNtrRRsxbwr7ipBFDaJY1pjGI6ArEDxtcW7el+EPtcBj443F6lPsbhjF
gd1yReZF3qo7cmAB66TXdFlewDEmtSgxzyhH2vArMNBqF7cJmPlrIVKLkeDDcYB+vr1QYRWJbkQK
6A7xcqa0Joiqp/rCEeya/SFrTe8S4WRZfjkDsKxmJeWLbQF1Fu/IxBsaCgogs81z5o+7Qf+SaRx9
X322JRbBnQIaVR/t5mrpvQcTx/CPCLaTTbaanCuWsJBPTScuk50OFiTRxTwR3e56pagXpRcONKB2
dqaD/jISuWDk/ov7iAm1mfXEciTrPXjOWD4J8r5OL7bg8ZivDH/gge1Uj/FnrtFcZkI1a0BBYlog
zovfLO2AsKe0iWo1RXChSCn1n0osULUGfWlMx4n9KPVYDdG5xIHPNbdrv2uWou7UQG+Bth0uHbmu
gxU7xvIsKHJTSML4cIpbZCUoPWG5J/+YdtIatGrn6bcnAdndClXNbTOkgDIaituIBxKTdQquDWJi
ZVna1U+3BUTTVmFj9K3LLZy5RN3b0DFvLgBi754HLtJU+wZqBNKwEI/ONv2y4wJdc1Gx/8kQa5zM
+tCrrf+6l7+LWWXlOaQaH/gVxZ+CVZP8Qcw3+Hyp4Vdm953o+dE/MuAe72Y63RLD21SM20XYpQbg
jLTugIm726eNjKSp4vaS3jcTF+eOzOCRk4yfIQmsBXUojabqfp4JPOBk58l8WwFZzWo0PkxPpvGJ
kRqpivSYzvPrCQDiG9zNyC/73L6+hoU+FQCXnw99+HOYw96JlzHqIJGEZKo7USwRIlTN4Ew04ZhX
co9o4TgD2IvyFSBi1QJbJix8XjMW0fSEgRCYr/sF4683rFe5x94ios5Dtxpc1J8SeIVsGgA1vB9Z
dXq3Z1MBusMuRlQ86YScRg900kUb0zvSWC0Ty92IhkE0Z/WTwdwdtS5pKUhUOXV4on8hn7DPujHE
Fi8yqjI3PYeSZdPWjwxgapxJ83+/0d6GOQsjWaaDYjPHRZSkOh2AUTFnFlQIRdCNb7MTLqQJpI/e
1rOnV//ItpRCaP3F5zbfysURklK2UpCi7n0w0Xiig9L8ee3FMU9TlL2kSnmfQjFaHe2gOBrnbszU
nowxtMZmNkJYDbWFYyVAYGTwHE13elFSUK9xuMMhdxDWP0qP2+0uwY+L5RaK1RBwcn8wYSHL20lX
sHMkc0XKGE1/QUEvF/lJMURAm19lLSFWEibb/bcYgena9iyDuicCNSG08fdi6aPT9mTqd0hy2L/0
3G8RPq7W/ivjDluzW/hcPCuJiQ8lvJsm+iv0N4aNmAa06KHLc7YvVxJREET45s2pEwoOKVL4gdrV
Ris3ROQcAP1iTwZwex7fN6X+IuZYtt9W2kmL4Db5h+XRsspRZJ48ppn/7SUmA4SLHXCUqGB9Ytr2
VHyLp2G1+yvAcw7heCv4UV1blizp7XOHiqZ4wdemv3Zgqni5EqdrRWuWYto8nhFxslv3UPicbeq0
EfhTKlXsgSmp43NGf8NJW/5VACSPyYVsrQ4Cf2J7RdwyzoJSq7k0tWAT6S6OTisuKvporxJioK4c
eq2FajyfJYrlsz4VyfdZ2eLOswigRVzU/mhsYM1zJfLoKEnfDzS7yC7GWbLqeqMJzaP9aG8IhvPG
DLJRB9Dn9xKHNiEQfgCk8EqM4RlnA3j9qhFL3wZ/ij/ZvtkAMb/1XacJbcWi/Gcklz2XfBrO89Ke
0h2W/fhLQUOTRLjj3SEPuB4yTxpwY1PllHSDTCCJGCaxMFEZ8ATd4rjzM9qNAGj+NDmXmje6Efad
ZaBKSD3XS909kckv2oW2ToevMxxcHyEKph8l7MA95VS+Z1nnKOeHPfZakHbrZbJlZojTXVAnbEK4
p89/TcGna4XrLntssNEXRdtxCdsvK0fPsavMeSkOD2WDXlb3GmwVmRzvWnLcfSD/ggOkDPAQ56hE
POEcS3Ya7c3W31TZTTCuk9qD2cNziCiV8+TuUiNyUN+QahVT8hTn6oqiAAtSVCuSFmo9BGUaPAC/
Xj909boPw1YhHO2YVKJYdD6gAj9A0IIB2AzsvH+Jr5ZUmzEjLSRHAwl2oENrYACgr4BmGC0HRWy8
fAGdrpVPiTKLnk76aOk3/wDdsjV5N0gylj4OiMSyVAaANaQMmn0It2f0b9umYBb+fsiBtvy0BPUd
misaUqg8aDrrxBbv+7BUVpTvDTjHABSsofxLYSscWBxjMuJIJkjb+/d7SR9FNLl4qF00+rc2vzdf
Us8POychpFc+wAAAbfv9M/TklHeqr1Byj3rlh6HYcbTWG5GIvH42Gq2H0GDQSUMdoPNRkrD9T5Hp
PxizgfhJDV+vxbEMD7NazD/L4ph0yYAgLcx99OOZF7QVv35xn6evKeI3GW543kTZYIGKpo2Ghwiy
DXJMqCJz9RXPxHN2JEKD2e5+wmuR5DLtRVZxVQ4Y3046ZFlXTF+7YNCQX+YLZeplYYqnYd4pT33k
E9u3eJPBUgzryYt+RoCs7rybn3qHTCYass1Q1KOeBBgadrvyWDL3RgV6nEm/fMEgrIpsZPrpbAym
FbF8PrglnIuDk/7KEMxHn1MCw5Q+J5r+d4llurY/Wr84aM4BRc7zo3vLlnWjugGYex8woyTXrDtV
PcjWpHtMNjOva/F7FZgqwPydpGWKvWKRYtS8XB38INKj1qsLRY8fAYbSujlSXfufTopiRuAzskeR
XYiJpbfoStzhjWMsXEcDroYgkV2EGcc/YLhmZQmVEfpWAEc0MZirwYZPmj1l5D+XRMalmLPpusc9
qo4pt8lmZqYyCcmk3kvA5K2JHHRhfMFDpa7q6uIE2DqfFBGNMGs0KFK/qtSVbXYJ38g+/fabh/Xw
WcwdReMQEjQL8HvcToNY2am6Fcl7+pXklpBUXLodT68CorDKA5e9YsvuoS47UF7TTNgO6XQ3mq2V
r8S0HrC+/mwoPbm8eW2kotxZreWxuH0bc9AU31aGjjkgclEtNY+0z+kXDRSvRS5y9XxnEubhu4PU
8glZAd3Weimt77+78tkYovNuvNNtI5rmtxZ3+oiXHEE9gYKEWDdpWthnaNyZ69zRBbJoqTvDnEdh
ALe1wQIdI5FhskLiGBCnADL9GB+kRSmzbTIqOoFIr7yEfYaisgjfBfIyWQAVlkJH0L0ouZd/c3W2
pHvuEbqE6t+JcaeqHT9EgPNuAlVMDJEpDCZzmhWlgwtfl/auNyyEjwlP0J0hBxz6Kc3jWEVXQufH
Mlxj6+NsZqGNWEs8+W0WruWB7Xt1gMAqlrSGLwceRoVm8L0Oh2ANnKhIl83QyPG0h5rYZ3ybu8GV
o4198fNpLPOL/D6MwsG1cmE8kDGF6y+J0NpdfJTTNDpuNtB/5tcjnxZmN4IN/OvB0vNgHcaSI1VX
CTQO3R8gqwUvpG3QXBsy5mMM6IRKXTx80KlQ98LjeF1PeKCF6rfrCtVIltvAE9QrV0K0AeEFO7r3
mDDdazA65b6Bwlrdrz1RcMTj1wiRllKxv722z0Wgdut6BjZlEaWFKIGitxldL7Qz12QGKcbfhiO8
st8VMKsZofJhYSLtYYr06xJH2scXPRCwGwEAKq3H7K6u9VSlT6HkKi8/xSub2ij8cj5dEYX4DN5n
/4WbaNdPeELZHKnTpdIne+DytoxJs0nY166BZCmc0wN6gy0uUGkCG+bw53LrdJ+ZXS7FWvKODq3W
Ud9QGtlwGsWvW9AsxqRW6ZtevMBn24IrMoJv6O+/F0yeu8Ej22xvUyGAPT6VQcyf1i0p5maqGMn/
lykkG3P4bqrOZCcMea39mI4kWroHB0OCO9+NF5Pv0Rq/mQQyoAuL/k4DRjSE7+tuIjuZe9kFKkgI
Gyqi/V+yxyQ8CXNTWVtgPxe94Ol9JuguuAD+q1eLghUprGPu7aV3PDmyCieubA2np9I7kWlxogha
sspDP38BimcghXr/aLwNyhF5oSvRdYioY2mmx0o2ZZ7orVyLn5cdqQXHtiX9BpgoWtAjyWZanbEw
kVKYxROYINs8k7PH/+zSVPE8iaA5UCdK+aK6x/+rmtJXlG63+wqv+DxlChclYRQlUfkHRMHxp3HK
xtNj6tl/S96omtXXOnFTsMpQOsrn1Wd1phKSKDAlnAcMVU9ye1NwBT6/1oj7DRY5xC697WAOTv1Q
SWX55XuVMOqAnV8DyZl9CHPecWNziYDn5Sfd1SwTNkzWFQdnLA74Y60g0r1tBcf/AWeSXHv+iUaD
r/G/KLrOBFk7KzN+7TrRtqE2RI59pywLrLUA5WgyyZx7+1RKy25WVGIKxjVSos5lCjEF1MhW6nau
wJ9eIv7RV1iJ3K8qJ+wJH6lTyC+bFOq9U8VlYTGEQiii7zLea3PRPXBue+JC23UX/CWpjGJfA9os
Ny3mqP30Tx14kNsGYy/OD1zOGUwaxmz85Fe5biP+IsJS4fhH/nOjgdSH7mENpT9u4ATSuk9CqU+n
vXKYvoOhGHptOzvNrBzJl+jtcDWtWgMemzR6DU8+4+8ruX8broFZGKhndgECcl+C97H2FKrDRGkG
XN7CoawKIoRSzoRiOpzJ0f1uAYIpQP9xIOCeyZx++pakNlRcWCf0no7n4lCe5272EjFQPVFFaEYR
b+YZnGM628aZdRe9HFUs5OitB3D5Z3j3OKGzSnjkYZnMRq6Fb7QgN/0Gz0YiC56fdDMHP2Up3Gut
U98FLytm2PKwwNftq48HtoIYQWMXvca4PVEEvreoQdnJ+j1g+OIc+OmbDx9F39oc20aA1c+pOkTC
m8zw+9HmJTiolizgGx0pjP10PzZll5aG+FLtPuoJb9rtsWlAwsgnRrcLOi0TRgOdXmjtacYrqyGJ
j07xC5UaL+cPR+ZtLQSqUXdEeNooDOcilHJyyZwIi3hGr7epYlz8ClGm1kPX+JO5CKMIQM5W2IUT
Owwf6QqH8pHtuKvJ9+abtY1X7Z+pYZ1Wm3OdXCI1gfZyvavUeFrycwIeI3Ola3VK56OiGo2jCmZj
SOCQ+lwPnYlzhpnr8I/3ooYIjtg8JTZDLOGsMp9HmtXYhbJzY6hHnhDXQUHlk6nbMqu/cXCQzYMl
unQ+iDsKlA7HYqRXw5Jne5C6DmYPE+vEpxNIjBy+wKJkmCf1R4o7JI8y0Noth41UrjiGED5HIEqb
Glxl2X4MCcZ7TcxiVe9sMlswlB7w0Z71VE0F7OmVc5ENAXKzDQSomlt2iEOK7GFd49O7b5joazCw
LBjMt0Z1h93ZjekW5dUU2SyG2WTGHx+CvkWevl6pgn28NUmmBK6Bv2NZP2PRpGlGz75XMFqBwESM
KOa66TcmOR55tIsz6nc4XfL7L+3i4CVIMeGZ87uAmWj2+lzvirAjbP75kOho9YyD2ngKZ6s7gVrS
D+jkJtGqsfXXweq4rFZH1lAz5ze44gyCNKQn+M1n68ZjBUnvMWjxtQpyv9zz2kxhqPMXiitPtdAJ
Eo5wkm2wldBfVRoKl/7GXHtp303hB2/RzZadF/yjxdCHn0BmTliI6FiJucuuIme0WztcjrFnybh0
E6VU7nYj/n8Vz23InYuBpUnVXd8x+xXEyjtqcwh5nXmtC0+oJP8Qlo4HsEuw2ZfmpYWTEh6VMJqN
dcRwMchm+s6F3YMwsE+gHCGhSQg/NQ7IGPcPxZtr5MZNPcGCUOlvebOIy9e+eespU0243H7HcvbJ
fX9qfTzY7s5spzzVZnCjObKm7ueyjATucWkOj9saclXFzUDjkuVEolYhqarmdtQy1Jpzl84VA53x
PTeUwHY+3X1WFWrxZqOGgM1Xf77wvVlBVyRTNSiOloCZaMmm9RHuKKFtRDow2AkMwKsdRb0Jja8C
qx1xIaQYvrOx9byKq3om2bUgcth5EpHtNrjF+QFQwwp1CfaUEWrPFL5nvQg0hVlPfoh/aKofuGI/
7GMoSHFcFcgukYXs4PpNAjzDFnA+5iKkPLchPvxKX2JaDOUr/VHUIudcQ2GfNXuAsCPZt3flwVRw
OPQJtsmtJXhzAKjV2PlBkj+ZW6Y9fz00R4WZka/o3mfYrl1HQJuxLN6BTGRsPouIw1oo6g+U/2WO
krAOo2/GdAUdwCPX3CIYar+xOkPoVUurepma8TjL4i3OJojYCYKHS0CinQlRI9ZkEm4g4nAUvWO9
qwxSh/CQjwfoIDu+qyupO/6nBp3S/NpDzpAxBws0OoOxmdnYVRg/poAweyFihkNG6+FBakFpTV9/
o3d4nm3AQXOl6xnAg2mkrosszjKnlWXXvKvzJNchOzAAclYRo4lg4D6deUr4X7OBUPXojGjlo/PT
oo54PP5FoC8oKDEpYrNZDorX+3j/44xaBIwD7BRZY2x0qtMu/mfYHxNdItKlx322z2TuyIVuV5oN
c8K4jjDuhV4c5G7JER6FtcRE3cDFGUZB1biuoX9k/vNlPBw50INm8ZC52N6HkChejbSqTWV9y5Bc
zDpJcuAagblPPwLknwDd+jd7rroPtPtTSeWbM6Skfj/jQxGs3WQBOXzolRbIRbSg+88Yp+bI3sd5
+Ps9ntGjAhqQZ5KOgNQYTWFZXul//DGy3cR1XZHkckx9to66eCgGq3jHLkK/wH+np5hez+Ytrv7N
Q3e2v8YVxY88eHEsnfbRI0XHWa+TcHxy3Zz+WqcZow0jOt/kmNCpYVGbLSjPkA9xtmePQHyvwq9D
BUdYB2Ft2PFRum2Jafc5R4cCCoW49kSikHoLY9krBMZJzShEhoItKLJrXuPY0QvOsxI0FfFNoffg
i0DW8AugGldUBnkxqHMMMrMhYqE6fza5/ChphNri4riQmK0T9R6S3bNcnNjJaJ7NRuNUTS0tKcse
t8MXMRLZ01XJY8ckwgtPki50iKBQbMUq/nKi+xbbXSfwf82L0a4t11yOcbbBnbwz5+6HElV0cXhW
DmKf53KUR/TCFS6T4C2GLKpkb66L+advxChAXdXYjhkxZoOBFIBBx9murqex9AS8VFuLWG1eUuDR
FC3TPx/AddqCJ8mgQpkXafhGXK/T0d+b9qHcX0CIpqiVlP4mhjpN5C3eMRY4VSw4BpGVqgB8CHdo
g2llDJt8vB9c5oNg6bP6c0mcvLuM4hd1a3TrX53fAwEsAiW/aqQwNE2+osoq1Hz98C1F7fAiYwjX
L8BFJ+8L9NHMrM18BV8gU6I8DnkzmPKs95hLj9wwnCK+B/6V0DExpidnFDr60t8XkdWQuJTPHRom
w2wUsDkJYzPztJcXghctQRPjStQVGHqOYVDhKyosWlBbCi4p4Ghob1CsHaSijnvnTCH9wfit4DFe
Sme9Zk3jQv51AHAUJuZYsDg7ayGo3leTF5BQLhPv+YbrwrFq8Om2HXqqBVYjNAR8JOdPqIxSewMN
+Qtu73mrIRKJxErsCPYpH7jEWvXotlONR7/3tKuuTJzfsvu7WivkhJpDdoHMaAu8L7nGf3N2GGQO
c/zC9eGJF540X00//5L/luFQC089hIShC/JLwlBbCwgpTP+QHK8BIxgeN3B+IiqKnOv7vnJmWe8w
bDJ51k4v7Uvfzn47l/m/nX8uqCGIV66qVtstA7jESa1kjopgV8SwIcSXr76mBSCuNbIYlTG3LI5o
9Pils4KQDQk6Cz4CR1AD/1YUkR6CKaf5Mz6ic2xPI3rTW33D60bmVrmwKnLo4genKAM3cH6Ytog4
goUb4ksz8/ovBbms0/P3JECgcfZRP7RDe2CjIozpZCH1XJqTLkcAK37qW/EzgTlQtOFC8dXr8pMj
waOBOjQlal2yeSB61RkU0SFwNyBpWyBWLXaKnB/s/823LtoRtElfHjIyL4QwEo7toTP0kiUx/G8L
YXz4Dk7GCwyWSNH0cR+nnVd4w2mGbyaXIlH/1VQaQmO+xzykZhV3fELZ0XAjP0DAQ5UYuawQZGoR
zwV5i5ixeL5ba/I1goV6m7WnzxG4dlB+Ig3qVBGy8QzCX3JkTjeZy/W2Md6RFEjwadf0eXDkv+eS
IeDQsMmwE7yUjHGsp09YC1pGaD3SkucAbkfdKtRrJI5meWXwTrMS2Y510yUl7oiIpHjaR4piDVWe
0mfwGdlJR7ElMzPQx78PwcDvA3PxY4StexTWIVq3tHzacVdIJjXyZvsl0SfoRxasg1+t7klgcc6V
wuy40HNVHgJCvRzvvCovo36A9qqdqHIKgjA0vVgo6cOfqs+1IK2dvogfzA2Z0p7TCxJqnvxRG9rN
1Td/2zmn9sN4Wrm0iAg34D6lO5+hC15EZsctFxJajv1DGMHSLCjeYwPtRFe4yKDeP/L08YacNg0C
sU63SZxoiuOB+ZjZk33WHZ5VTK6Gp0QsyepFKTzkcE8k0Yk68jmngGOb+YE8JFu5ldirsll5k1xv
8cKogQDuo71l7YqGTmU5OnHPF7rJBEvxOhQ/NdClcxSkVSG1YTkNyH+6Kn/WTctlM/4KmOKy5Tdc
6RN4Ad9W7JOhC8hYhvMSDYYZRIPE3/hOL0AG4WZsAZ3DkKA4soxkt9R3FQmxA7xu03PdP5+la/CT
xIEiqfe1kHjuhrM94+ADkn6M53O+ATm5SzIh54rfmTMqzVqxwtQFJXOEA2OB2SooIqhdY4XrluVj
TfF/eZM8pqM5eZ83BNaMciCNo7YTQqZG3RJ7dwUOJZCnDoqZpQgT/SPTlmebk4XaoAMJWpX4csRT
xi32SJNi+MQuQvvXgiQvvEE4lwx5XjZJlvBeH1/EKcqMJCVu/iksFC1UFvOE5S3s+PkJ0Egl46CT
arLg/QNZv1mD0iYyTcB+LUkJgTAw6LsQ53WC98/GqNht6ZVxRkRJWsG1ybGQpcIUuiVCEPxBjPKN
8HP+2vj9L1gkvBXgODEUaHlVJLSziYAi8QmkWQDRUUJRkrio3bZnhF18JM11mpRwIkDGAplqJOK4
4bcSsbL+r8YgNbob0GM5GvvrBKAEsjncqe1bsEwLAyxf8oQz2mIOHFqyudnzVDR2U64YI9Enn+ah
q6YUOgGC0LswhuEyznBDqA6dE/87U27t5STkhT4XtNggSo1AjEPQEyMCSwcdlycLPZB4y/wSYYdZ
Ood+B9e8TtwNtt4MT/dOnviCb2pUuqsI9EN9GmA0ir3CShXHRu/14VFuHQzjJSwQ+r2InrwUC1LP
Hb2XXOuKzj/XV3brwYjzBJm1J5CfoGJpY+LDnOc4NG4GYOp6TxZparaCuPLNL0qCTl090ebpnjU1
LgeGN7+QNXdjtFdXk7OnZ58MtdfGPAJoK8nMvjHdhC4s6qaOuGB0ks3zFQg82V/vKm3L1v1nRTiY
QajY0U93PGEM+cffmrafH8eEq6pMqA9Osu+mFEHI7oFsIaay6oYdbDReZnVJeAduZXQu6KkNQNgU
yKbeR1catI3rFWcQvC1Nd2abEv8qdzS1m8jEJHF1+O4lPxP4exGWwxGqxBIh4lW2hNATWZT1O4I0
Bl4TBrY0plg3BNHAwicAe/J7JK+1vOhnI9aHfZgeWH4R4UA+/L9Fo8XZ58b/inH/i8czErF4o9Yg
J1si5L6wT0bBmE1XEn+8Z+/5ZweReEy2+BjchxZwJjUi9+rBTWUluCnfQRFZNdCFCru254GExMks
OoGpeTxWvQQ7hB9E12ya7mryF3OjolsOTYumBcv0OPR8i2SVH+LPXOv+dQovMhuEW93ZLPkwhSxF
wNPL/7OmWnUBD1jzoQT6QS0QW/fRgTDsgySzvA+OWGsdKpvKKBUnG2J946kuxA7KR5HDYnX7L1ZK
7bH+d3W9xHtwXfOXRc1ofyXUpYbVhiJgSZ1VajEnEK+CW4yo6Ci+XebDYkZN8Wo8vELC3HPpZJKF
BQ23BliWU0qHAJF8WufHpahRrAXbdadWq4gc/mORK6K+E34W8QsnHcJ+sUYBaqaqmeSBMEl4aufk
f0qwkUEtQaVasasTo6XAnSw6vGXPSaSae97DGire6my3H72fj4EG0T5xwMab00dg95YLj6SeoRuK
nOMYoYQ05MTe/ej/kPSXiBH1bWlev3XiZhIIWHPm29mf1CCbS2z3HqeVtrKBnDAjvqTdL8Uez2me
BdI1EtryEuVcf5y4kTVyrRm3l3PcNHntRHNBirxeQZfJjJAmXibNcYJnq9Q8OEOHp0yyErcxl/rF
6GMGEW8OsN3rcwqtkZJ03NjY2OIeBLLc93VG0cTJOz4UG8DvHsnn5H2bkQuxLEhU6u5+IWX6VVMR
zhS8pxj0IHcARPfsEp+5ESQy5Ia/LPGFLwWWmaq72UD65j+rc/ytgwDDNhCiT9Ka9eNjlDK08GbS
sQn6E5m+6rzH3jn0OGjzB7XlxJmEUXykbCqBmgHen81E0xvw71WxcbdBgGssyFP+tpGF5242X0Zx
0AeWUM+VI3qFVU9eOlxS2qCRfxf3SY5nZydBx9mWeRDLCyaoSDTUFjB7g0kuLQ9sER4QW0+KU4ub
UiBp1B5lZaWykb0245pIGIAxZDciZLwoJs42bddNkl9xlehunVJZQyZpwQlX2hbnQK6w1iBc2g4B
IC1e+P/bhaUrqHyvJO44dTtnCKGRuzRuig90iZ9crQ3NnrDYu/WdoEbDp2OPLrsqvY7LUdcpV7zL
zxImN5fMo+TuKdR65iS2T3qrNz/qFi1xLHrGfdXWkuoAEGT7vIjQg/Ldd90Dcn/FXrI+TxEGMYLo
1ejcT4Fc5uI6QFhUdSzfenK4fskeYvH+J8523sb5G4KH8B/C0x2opTXrCd4X/6ZjMblezBL396/d
3/1RY9LGCuBI74dK4LAvbgYGFxY0bjwoWJyxe+iArhjY2/UcuiX1wv7CbLuXXg56vhvlv/CVomqK
LldSHqiFETChNCbX6PfvkAa7uKyxCoirvjnO82YR3vVoyKzYoSUpuXQyXT8SuD1R8CO7xhY+P3xY
if2ok2cuXusijRR7KlSfG58gFQDr94d5xktpzG5lnJVh42S8l0Tnbptj3wo6Wy0Dv5vejPkrYyUR
aJ+sU6vY7TplsPDVqQUwD5g+tx3fiZCAQ/wr78OmMzgM5M585K+8eeT2i4Xy4YVlT62E0MyHn4WO
/q73EDMMQ33a3y0roCbYg1TFQaBDQ/JGVLHfe7qNfOzIrvuUTH1ktTaf4ZhBRd8Av3HQDSNiT0BZ
tRBA5Mm0b0zuty8EvJjp5pcoPKYuE/HbnIBb4QtJrzikMWI1SnnBD3eBq19nTitmXA7+YlrgKdWa
jcHXCgzMz6KVglHP8823fQWeRh2U9+IdT+6xsjRejvTOCaBDBi8cldtIBLori1osZz8vmpBajUFt
HwZhTPcr8cJuTQYYNVoBQvYrVq6nAvEMpcqTQBl7DwKjcj3eRS8gvNdDct0jE1+G4MiayXAf4n8O
9AEoViAm5jCnTcMDxR406FmqLd4q8LsRyh1IuVQPGXe5ABl37AU4zpQL7+ReCs9+kM3D9wtsakhh
b1ZZfigT2BpGHHeSmxg4XNIjfBcjDDcMx/cQvZO9W0wwdHEqnjCzyP6tMoJ8CN9PgXoF01Us6l0M
opkWgkoDth+g7ftRkCt+VN0+Rm50vGO7xnoA9oeXXFUMXjJG/QNPxI43c7Ak9oC4iP/1all+8uqo
GH8717sklI0xkuHR3OcIynqlhyCHbQcSSNQ0fL4lc1Ab9mu+CzC0+8bxobD1pXiOmzrtv5HtIiAf
dooB6DKElK4VivXGxk/Yo7lqzW7UxLGvZUKU6D2Zx9WsW7tQNUAbBvYe+d1Q/EFGjL42lKmJ0PFj
PVrktstTgYWvd8yAZFqHw5RCXLaimEFk7x7wCZQ0wb63tEV6w5jY79kMj1SEZaMCTMH7pHSzJpfU
46KURPxZf5KBr5Sl/w9xacWIpTD7tg0AxvD0UsjKAHQKUoHjsXHSyQZLCxcjqQm1VvRIMon89Jlk
0zxWxq9P2wfa4bL8vEqO6XDX/YoNrH0IjGLaezWOApbZviF9AECQj1pdTXqv62mV7QV0YVd1uLID
juqAp0cco20tQa0EoWuWkGy3JSUoYKpkYWh8ecSsQGlr8tzFWmH/ro0f/1xbACMnuxDWrOrRfWfT
seB3g7tAzhtPxma24VtITqSAmkxrTI8r01DdQYPRjuWjJWZsNFX5DsBjCaHBON+qS1w6/Wi6wD7L
sKTmifctDiOZecqZfLjOxJkRmDnTo5kf3uyd+YMmZlSMzZLdRtDX01eOtuozdaVfZapjthJ8/D2r
3S3w+aI1T4NMWqx2ljxC1eU8Qtv0PLHs7UMsTMst5BQ6i7b2LVzG09ZeQ4WNSTReRWwX+KyjR0ip
Iqc7Zeh3Y6aLezJ8rRJKQMOUEwSl+yjm2qmSH+lSmGZphIh6Jvwv8tkLbVb3huLRuI+P81jvrl+m
RoUecWqNqu5ZSA1bGN5hHC3+BBOxfZUcaFlD4NW6SzC++aVbzVIAi7MMuHoVEd4C20TW3SlHLebd
ezzJYRXNIeYnJmpwRttJq26IJD36T5R1asjYRuCcVSKMLclZklrv/Ec+24l/mC1WGypNOD4cdWe1
B/g08MnRQkgOAnXHQNI+/np/2cmpez3sXBmCndjH4GHx5i5er5H49d/+bduuRBBczyfssjrsVLOR
eXiytNm00vpku7JVU82DoYGFVRtf1pdLXCw3yaZhrzDHM7Q3rwaZuNmWnLgJq5oKDXzZfzOCTyOD
7ueLe8OnkFSfcS6X3FJiCNOdqdlMj22UhvBhBjPr/BJ5oNq/2s8pWoad994RVrSIiQUDXzJNh5Ql
sAB96mE6I7uTz4SuE/iwjzT7AA/s4ghigIFFdHpuTIPNZ39NBjMbw+opbgKfF0xH69wfntIU08ME
mXrng7zKG7LPWL4E7E5oSE4eLu0uJyy0hOtSXTqsRaaam2o6EFhsJh2hX1XbP3IpWAduVoJitmk9
GvuhFvnlEvlnTDXrLQhRsnw5yNSNJcMa42gOBrt07UQ/smKohCv7J1ixMzjdniLviAanb4U6IqoE
0OCoXFT+utulAL1OkiZDoLaOy58ZEg4ZHzE3o0UOopzlrwuEvAEbAhd9IUS94qe0+7VIgHRtmcSF
Q27ATJk3NAmIzRpYgeXLmoU4hqsk4BdA1UtewGT/pDKGRCmHNtCuLKMIUMgkDslRxzIMjyPlxinQ
cufNDdkVllGHGKBJxPi55VxrpcGT82S+ec50k9Ggbdn/3q5vSnR0sENveyaAKpaxjXqDKew/Zrnw
VFkRaedaD7TFgfHcLfbTvrRlWcHSzmGhVr7hNqKa/bYsDP+PbGxIUSeI44m8a6REFI8onCnezRmh
J9p0BrkbZn5F0u2ueVP4CSvBxy9IDhgxdeu2wE106cegn2IPfVrnU3xMUl9TSEcm/IKWvRQKDQ0Q
HNJOHY65x2VxfbJYawKaQajf78j+ddQ9rgmyLsOBMLT9/7+Jk/r6K0PYQKKwzIlgDyFxsZIifsuS
PxjE4FWdnjvNQeMgVDBBw9O4KfZW4+XtsNCo+05/Vw9XLZQDC5YvHdS0ErMLC4xyAZa55/qwDaCb
FYaiQAYsyVad2fBrrG7kR8YiqCLIz7w/dUr6RTHjufSJZUmIr+B9oiALaQajek3GiXmQjByoGgU/
Yd7V2T+z8TBGvW1/4MUlD/49b7OpJqM+kcjpoDMtEj7k7Jg4MTL852xtwvCB7i3FsfFdoAtdnEzM
0Edr4vcYJU1QM2f6wAnuTV4JdA3+w7XnxFJWcpGgqlks5eHzF0yS5i8TIrvO2Vz39qrTZ6EFyvoD
BqfyHauw3sZ6GnAlJd+J5FKpjJC7dHRaaT9IiAh9jkBUpqMLKXfNB0fBc5Prsu73SnwGXiblcCJf
if/h+nQUrlGygpO3m4clTcJTyLjq2SNnpJ8Q3Ih/NDJ8aWnOkkt88RuvXZEjqshxZjQNib8vkw+y
8Co11ttxLaoWFSDNqniOQsvqTKASXDqYvj7lxLgJN4VzsUqurTNnGyoWC/N+5GB8+wyNA8Hx3HrM
QASZ2KsDKcwBXeaoyZ3/F0kv3amBhVn01kByjZhLfxXhGcx7srQhtdpATD1P4xcrvB7ATe7d+H5/
eL6TOgByg85Uv2W4EmJDU9DVOm27Mp3bSXRIIErjkcTi76qhgwVdzqVoXcxLB7w87Uxy+SQ4LWPr
SoS1Wec2pn/1jIqrtQIS1r4sqvXh4725pe/+uKpcFiGMOKyJu13VeP8JIgYS01WDB9rT6eXf02O2
LuDOawJGr/FfD3YfW3hoDTtzjRcL7R3wyL89WoBsKhBfSXsLYRc2QIAba7n8pBcltz5XDB+BDDhr
CNXFFZg78vv5/CHsyZpuNBEk0aQEgnjA+gtIeYN8orWjDoJ54pATF4ecyT8OxH883DXI63YtD3TL
SB/xpnSO2VMqHPhs5c+ZZHsiHQRbqxC1dGfwfoJgE++Wx9h+nesW5kQkd52HFVl36fpOCYrm5iBS
e3eQvoi40Z0PTebw1+pbbAOl4XIfGERtsMZ8Gz+UC5n+vKpL4YUEe9JQ7+oQ4/Aym48yd9dZyPP7
FTxVnV6tV/KXI9UVdFaY+SGP95UzgQgq4FwvSjWMuXex40JqKIgrI4XngstCAY3pGKOoetNIEINr
9ruV9TGgiPbdHb2owhlmYybynclPQzMxeDyAR3qQ7aQWhlZfqDNEqGRPa90agP/Z7j2MR4of5Off
eRwQlw881oGZh+Jl0C7WStV6BuH49rmMRe/H/XreB+hrOC1xuo9u8AwLG+DFOhWBnJKhGgGKjKN5
CuW8tmwMxJK7sxD5AXXA0417qLYsi3t89TA+D+coD7WtkSeUMiAXwpJuYVG74WReDavgxiqdNnzw
xE8uLEWod4AY16dxfDW0rq24iPxGF0gWLEsIcs6F2g2wR4xdcUZnr6NaFPFyzdtATuN9HzNVXcMk
iOfLlYznIt8TFyCamD2k05+TrjsiOGdmWJcuAcx5SWAMBQcylUqAiJMvJajL96DsOktTkIiAkpZU
XP4KrAlGi7nIL2eC784xAKdopcPTz5F4HihyCNni0hBGN5LMgAYTrFl53ju27hM9uZ/CBxer6FdW
iHwsxFW2MomCvXcQHumjLpbXrJ2rWSXIyJXr/Ttw4a++RUMI74lJcQAyqaGuuUQjzY6vE+RrCyzU
2Qy+XwPyrWfNYNJLcbIN4/0cTov0KVkKkzNZaPrqFazT32JYG9AyT3MhSU1gZ81/1KKy9gv68X97
Kc97KlMALricsjDGQ0erlMzktb03BtzH/KhdLo1Exu4pzJyaIsH6yqmt3ED9acK9+yGqkgIaUjrU
KeMGMQFCBjd3ddiq38Q3JFbWvwrFJDPvj3t+IVXj4O3xmTrYJ51yPl0ouxBEHAYv0mHFu/sxV7/2
UQc4+tqvT21gWYgHP5yVOawwOfi5u7zTvOpq19BNH6n8nwH/4d1QPK8i11HtEOtnj5FHWctpGS3s
lO/6abc0PVPAuZGkDvAML2PRoeoztYUyrleDwj8aHFxwZaCK5siNQRu+pNAZYBz2etM0Y6evBmvq
BmBCgEpCwjj8RcyaoNq5DvKBtKmPEEvzju5FSu6uG9aN2aXF6JOh6/k6vF52TyrPjnH5p5hQim8F
xs8F+ZJhNwxGIPRV/jYmXOIStngrzL/1Yb6NDqfKn+NsIkcSwnFbaX2e4RFr8+/FYeRE+PNGm+X3
6vnkoWB0xCzChuBWwPtokl6Ng5wYW4J5P2n5/UiKGW2o5Q+Wb7C/d9GxSz4HBgjcwpDxluB9wCBD
ADOWADuQGyqRXn8idPPtI/pYWXL6ZkMRxFOMNStZhEooAbtp7CGnAzKoal7nRexDWAhVxL8KnmQH
DM5d01BKAxRrYPWvwkFSyUzmkIzTqwwObZHevj3Y2Nlp+MJaidEbiCuRUM+Af+tYZqKp1t6z4AlI
jK6zCEXnf3TyjweuNrMJu+5buKV6smZUIRtC8HjJGAG9Quga7iBj6NFTi3Vm3XBRojy4+vlwk8sw
GTMUGT70TF/Gk+xKPCb1gtxpsG/3z/jDRU0PJ1OZRj44rXpLoVvLFkBZvyIs1IoFVD5Rn5h469Kb
rZlRFu29P4aKdqmtq9JaRKJzx1Cxnk+pCanxDi8iObPPQQLciTXY7/T9Q4Hp5EJY6yMf6AQWwvCq
qGA3vtCvP+85DJ9CwtkjEoEh3ZL2amtoQX8ns8UdzjgsERupVBYx/KIMUwZsoIA4x0LHCN4Jn7S1
jIJ8JyHheod2p9/6iJ20AbfFmeYoRj+vgwev2zOvZC+pP10j5flkzKkqcH02BXP+JFlsSbCdsASz
oJ+uvVEv/MSI4w0nWf90CpJ5LUuSV1Oc9jAIpP7fe3NI4/biQp4jsfdakpPFcdS7EtojyEK9C0ez
r5YWMNG3P18n98JeS2azu0M/SKthZ0Iz5akJzZuVaH4qiRbHXY0JHOhw+rGbR8D/mcAYdrvcEcRt
rRDlOag+Sarin52yCCLSGFEjuSFKRv0KZNks1IBEVUZFEacugTQTdqpG9qXcenskcCWSQr4IETu/
Bf692b923snNNO67wMwpwaFaMxMh6jGLHMf+iJXKbg/8w903q4zRRcDNOiVfmhMYwzb5zi5w5nQw
O0Fjn8K6TQ4Zn7Guqqfbu2nt+H+5HfM0lkSkoCwhZm3dlsxwdjV0wNxV4XbUmTOvCULMzkzi89LI
TkqK1Xh3nf4PdSCiGQZHBILYbXMNZ0a9F3cPt3pnLtUX6cEqMs0TgFGHSl5ZIT0XTYnKdSMw2xdg
nvJrzL5uw9Fs/YfIPjl63iZs/ZjVrIF8iS1CHwenBGHj2NddvCRpc5vCEJJntYPXUTsf+B3JWdDz
k+5OEFMqDaLxP3765D5MgBXX/0mIOBKxGMW6uuMxTUoH7pdwWP5MAFN/E9/Jjo31XLFAKyWTSvRP
junUPh4rIevfOXEDmn3qRpM4CkgGZBHtp1zLiHUraorcyvUaLOoc6XtMyOzghstB3gBgSPJhzySt
Ojee7RxDvAfhMjwM+oFABkMAzsBiikVb2EicCgui2JEf/bxTMWHYchTS3F7lgoPHaCPi/vjLqqdX
lRhjtokeBwt+pIKMNToNQiRojbV20aYqkijR6bIUVsAx72CICp++8VJ4p9OUDInuUycI63EYQ7hF
gnUGLW2VvzOHZdCPHCjTosz6OuBYoZIMzpQosjkQVucupxpXz5XUNYgJVmgmXA3NiXcc1DykUfBE
UkcS7n5WUkVWhf2cPu4l5nMk46Qsbc2c33N2WNLwuMPXeS3DGTJ61N0NH9qYJyqi2SfA+5F86K6M
UOGWf/mh6OQvPG4I6+kAZ7LoktNt1gNs8s44g95waM+nZXbVI8iaz6wVnN+eM2CvZysmDB7HNPZG
roenlochC3RPxQojuM6xKg0yBLm8fyO+CsOtG9bV+LtPQguk/zx0JBOuSPQyhPqLAyAKecSpgJ19
zA5+dAi0abIZb37VUPkX1OeTvDax1aOawKqcmW/BZVN/iCpIKq3rVGfG5TUcUDN8Au6wSYHuvxW0
vKqCZ6R8n2b+fmVy3wTayaO6b665YIK4MSnXkjVc0AYPL/Rb1XpEa+coj1WRQABFJli0g/Aw8utT
2Sh3KTgzSkTKwe2gLEKLc/csktd0JopdzzIG5EFDDw9zKCx9sRmAx63k6XeFrmg6J7wbafSkXQHr
VAwk8ce/fsXx35dtuT052z7iJrkCQKSGELHIoppK6IvDqxoOrTsqIbrpxTF+BnBGZlsoWfQxO7yV
Khx4tKMjCJ7kF4j+MtD7AQvxE4S2Twovy5xw0bL3thSsbz6wneJO0nY+cwe/wzaXFzAtUjMAwIb9
ftnV4pYCUEoJbHDuRWNXNqrlbXExgBfyKxZCKXLjbf9V80zdVt3FShJOCuRZ1waQP4/ukQVmw5Ah
xtsU3fb7Si1eU+s57rkFd2ZNv/qVLQA2xdNDu1jzyrWyeZIE6D/u9YHuYb9YUsLzYh9sMJG8nNKR
XKp2oX5tJSE255xjSqnmfsQqu4BNOIYgoV1tc9t5s1hLURoZvgewk/1uYLk8A17iKM0pWRWTF2IX
XiWk5CEkvMjGUM3+liwKin/2WwkfNhgIYfP3ouOy16/A+Lh99wRXPGqIO3FBuuqF+Ek7llBJLUM+
qu1Qsq76HgPI/K72yxy0og2QWB2QSIWKHkF0oPujjF78pYJs3LguqktG/Us9eEjrn7v1GEEaMdqu
CsEKxylKfXrv1djh47VxujooNrMxzU3D7gQNxZCLYZHKRnrRQt/Zw3HKRAIaSs8sfaXh6TzZvUQU
Pl29M1H+DBBgzrXpv/fv7Cw+Nq11CMoRW/RuHa7dZ3KfFQglknUBStFqiMlLh2KdrletQOPCBmFz
K17bNxRYcTu8VRMLhCqswVTdkM7LAyTBrDak1N/G2flKdTDasuShihV8eGmDkb6Vo9lD8ymgUT5R
TW9Sa28vzwPIEeO971cWxKomEjCM3oVY5rmRj2tmq5gLsvNL99g0NXzB4t1KxAC2uREp39L+JfS/
2C/VULHE4CxHk9npV3JvANN1cuvi8nNNd8WDb8PXqOQJNqJCuhThSiPMLXq5zfjmM7qbIIP6YJqJ
pl1ozOvNCN6OSHG3futAYP+J/84NWP19rciE6Klcc/OiQ183VVHe1jk+Ik7dhIClpTczZmdo0p3C
dlxl0rvFZaJYoYDcUWrFF8FqDMq4cg9vweszuStLaW3sn8ssxGgmrAkQTAWJYqJa5jbjF4ysEykc
WnhYVUd4A75/5nQWss8lPtKt7o79ALlaoCWf4FNflGmPG+FczH6+9Rhr/42UMrILt5lyWkVEOAJf
fbI5fD1GNFnaNZhpcSUfaW/5TyI4NLFL+n9ZhXPQ3nGU2pW4r4Fly/b28luAfZYqnPyrk4/GtT8M
2B9xjpVL/zJgzwyDFNy+yH+iV+UqtA3krtBq4xUpLt0D3nPyYDI6vIuTkAXP26H3l97MOPy0KYMN
C5sJ5mfA45i0Xk39kvTnCUEfHmCxxc0Koq1d4mx4E9yPEA6C7u6gJP1/N8le1aMfzGD0hAL0ckHP
IRQBSVQPHEH+zyvYSz+NtIwu66NdXEIrvF8K/ZtFEp6bUS0PVaoC4L0R3kkBXvulIoJKkE9dUozl
zh7t2jyHNwS8Z7KzGGowr0zwkm1oYaqskBeBbRChtHzZa6k8CNN2EVYM1BWlNJ85k9S9ZXpk1sGH
XvIpM9s219TV4nTUD+V1kqFoyFPj6MEisN3WoKRLYjNKIRY4bEKnHRouJUlyvYCfr9At05v3bCfd
rbB/s8XFfBXy7AfrZRdiVaixOJaQc9daZLvA6dhFdXEzlFzH1/3UuGG0qdOOtTV+tx8k2PX0ilZr
ETMFNoC9+UKS3PU3brLtEYvLUSkj7jbhpkyQMvOX4fL9/hGhxZUPcusLRw0RaZFtoLIcOwMPn2hc
81okedcxZu0AwzbhJu5rZHjyhJjr157GDplW/gcH4G/2XyBDMxNRCEicSa+3Ono3bUZgRmQ+I//s
axlMdjuipqaKjpMxOK3aBXSYzImc645nArqbjVrKmT6wfoCH++vDKqUBWWL8sFJS3aZk9D9IGbUF
fQsBVYMDB0oqtybiIszhQEJGTOeEzmFcWmBxoO0+62u2KX7X/cbHCLKVLQroIEFbKVF4Ri4ywd24
3ybSQvwq91nqE7t6Sd15oc+E7loLqziXXNNXlvBiHY2NzhBN7Ry8SQQbJ3g3ukyB6yD3QBBytTM6
U+LKhTROzz3UJH4YDXNWsdr6y5KqvDezBrRSjOL/DGB3N3QDYU5ofCPuuQKT5jk7te0sE/TnqZmY
wqvpuCal8W8TC5e3DsJRYGNS211Rw0HvDiPecFsIlkK3v0qAtDD38WjO266mYT9HCr5NKW+sDB16
e4cbmqzUpwbje0xT31XMf2aaCM1ehhu8QtEjBkzqnIlwM/F3SENIuldwTmf4as1d9Dbq8vLkNE7c
QTC6pacBeHcDSUZPXWea3qijwY7wF9sHQ4z/ArrEqLzv0KESKtG+zVOrGXWvl91l2CI4tMoc1gbc
ulI1C/soedffikPINmUI2ELfE5v0Tk6U04suFt40dYUAuZT3g3TPmHME9WlDyZtrmKOnoN6tbfB6
2gotLPZAmjLK4JK91xiq5Lqscy111chnTvDC1dP25wNcleLXZrP6+UwlW2kMDy/GEiuFrIWmF7aJ
Voch4xXMBNh0djHROV+xKAn6Ofqibozs9bjPEcLUykp3DekMFW3B4XEIxHu25FXkSujbKktAcZ1W
03zD6S1Rv59cYr7pvWUzzr9COZDMILizKlCn/gkJZknDXfY0rURf5+kd5uk/s++ym9/lRTK+EprG
mHbp13IrB6KxCjKedo2wI2XM7WQQEy/pPLWDUmFM80x9v0KfnYpcjaoyRGUgSyOrYC/IVTX8T//D
UV7w0Y+A6C9jQBNOtopZWFlqd+BTdtVbcEEAHJJkGVS+yXw/QaZtV7wp+OOU2wq/GsFcb+3PGyxr
+BhjwWoA6zwO4sXrsupTixlzTFIp77+6DqhndPrvENwO2fOCsHeaCyIEYFPZMs6g2CJO8XuhcV9K
CI2e1CxptTOos5exidfoRm7Y62VRjApTMiLIaairbqcCXHFzcYHQDb57BRX+lT3IXuowK0pYeQDx
eroq87Z/vJk/5B/VYL+RpEhJQTkr2kFBMiTWg2dbdmpUtezBEUIlU5EgegJqQY8bl0mcAKCis5pb
CeWvYXR97Sfj9aNEcKmgHrw0VvXkJ6Q9UA4zlY8tGxvTDP5v+fSTCpM81QreBKl0TuBqHiu/1jEl
FZAArtlvRyy/Vba/aivUK/Z5kqYUDla7aqvhgGwz9E34eX3dkQ+VsfBgfKVg5WiNpJjbdO0ZJ1Zg
i8cT23R2HWVZgRlDCcNl5+NkpYslfiSX+nupNuaARdzMB+UWVAq7335i2nR6I52LhSj0XA1wrqQF
jPz14F08GGYeXKu0VgDxXDlhHhbDoA69RBgI/7ezZr/PJV2TNwPyw7NAaW+R1DmRrwwRk2zcL4eB
mPaWEYY4fcEFzdoz2BYkqo6wVo0XkdPFimfvqu13s2mYKeZbMwb9iDe3hsj3XAN7FNF79BB8m+pN
yA4YWqG66Lc14ozNV7V774tPbTx3adtBYXejAQBnM8rpwsw1SYVEbPh7AxMe9YLstiu0BDbvEzQ6
eThZwBr6o6BtgCVmcesZ+hRq9lm/EJTNsuFPHU7eeyokk75M0Q+hH/HEgIH/JQj9UmEfSflwNIZd
zqYogJytzIECmAzkQftOCGWVQp9iWGhbnK6atfjIfrEdQnlhgMEErkTY3LTKfdqysFJXQxjIzGzq
GIP11RybegwaNs29bXFnPbU48xrTPPzPf/kN7Riod7Hh0A7O65d9dp6M6dVT65WdGyeJtlW1jG3g
sjT6ysYO3EoShHD3km0e9nt7mv6T18ZBSoMIUwEJd/iLZ6jcY7GQV0UKLzq/UAmZ4+1IbMsQT4i6
eBedNCTxo50YEhqJe0VaV3EJ2H8kSod1SHmGCYGGQiSmoFK/Qj4/USHMQ3Z7+XcbvkCP2V9SRLqi
yGEKlEQbG6z6B/xGWf08Wx4QnJFQlx+8rs6gJNjGsvEn8xJ3xfqmNXSYAUfhUkMSVo+DHnBubPjO
fkgqd3n/yWpyCUvyPZd3QILi86UZ2HPBd66wcq/VU5ivYyshJzORTSkIM46o0RV+bsrGUFaVaPfu
/2AmrkaAqMCvc0dPZY3KnPx3yBQVfiDitdu/zkrMPtCQW6VpwsPshZrwpWmGS8KFn1qEjwfql6B9
r49ZaYhRsiVPR+6DecFEoNeeYuj5rmu8GP+RIszioiG6d4d/LMAy2URdND8DrA4xeg1i5uHn1FPO
J8S/OHByYc+puS1UM+WUW6bVgFOXeWTaJhtiW89f8ahQ//NwYmh0LxyrrRJcDE+Te9sr1V+uljup
l6VAnpvJ6DFFg5rg1l31oFnhWNHq5QtNsInOqp6xbAPdS4iWCYlRcf8Uaz4Krccf1bCBt8cR1dxG
B8IKw8FgvFCkmmsL/K1z4bcbSVQbR4fS+8xrHQXziTBaR7ceq27NFRYo9ZTVGVen2XeaPibmzPbD
PJGQ7HEatXYsCu60TLnslHVuigkrQVY6iiz8jxSJ8RJzh11h/Y3m7g9g8QkwqcQfJbTLPECQjhWR
6s9C6aNo6TVNua5rt+ubgIBM65P9wJMzV46PCysXWGaDcJ9dVYGRq0D1WGL6NVgRBDPq7zdx17aR
OaEAvLzrGyIucG8dPSMJf17Hops+SksqL9+23Ei+0IA1i2TbDqiIYdG0KFQO4AB1d97g/RNE4/Fu
aGciUrz9c9Y4k7JRx2y7C3tMIUctzPnqv/R8YDdqfmLCE0p8fx6jY/+nETm5EoPmzUV/TSj/6MhR
TKPrGyLlCaPAvpscjsot9JOgIriaG7zNDH3VeE8SQ3aZ2dqxxEqtnw+noyq5ml0RCrzThG7rguQ/
OUjbebHg/85O2TuvWW6Z1zxUoC1wHeB2mZRoY5QUtW7LiROIYhqAVQdTre/B2dn325+JADdCDEtA
vCKoeoUREgCpZrp+zghFaDVzrULGo5lx3l48QAC1cuWGVSK2RroZN71HGWixW305NQl273+Az0JK
cnOcRk/c7NAI/FD7AkzTq1dl8CxkLWc+HVidZQd7Dz3mr/ehrfTuxNvUTJXiIhtnCcX/EmQTOst6
X92vsVL12YOeZoDW49c5c0Hr8sIitshR1zXiCthBlTQH7f+WkWrig3wkUvXUcotZthudDaGo2b3H
m7wID+vi+julqvpIwfPdtlDduvYt+rPuiSMtiOga3j6O4C6V7WV+hZLZT155faLs+SI6AQ251KP2
ecxD8Ze20RetjHKb3WjRlxEDA+0fZBl19NsW5uWRf/TW6hVxEq1dU6b1HAgYlDBD75t8KJH63gPl
MnMnN0Wh2IKB3TEwl68E3TxUGlqycaUNAfj6Vs1iJZHrjgQyukbb5r5PWgodjrQJW2IZvmG0JNYL
HhnKEtnExB7v+HYBpg3HaimxqlfrAenKMaDixC+vINOV9Y5PahKp51RgcRZ38CtJRp2ZB73FIAOS
bc3Ie0FTHURnOQSbV3Wnjh3YUcjn5gsfxUvm841nw+R98zEDKBDdu/q4ZL8e/5MfNuYHlWFRAXp7
vo8cWpS9RRVMAPdCT6xt8n3JkCr4QRzG2O1qQF8KojE9N74aQD+3ADvusT/mnRzHRVPnlJHYxPgf
QEJkH5aobOet6jzVM4b1wLhMC8W73acn3nL3EMy4fDs9hGUbH/gGBVrM75HjD2fKWIx/t+JcJwPL
bgPFmZdQ35sCObj+PSv2SHIrgmYmsjlWuApRl7wowEUHvEILtOHphlDsPsMdSuTlPwi3x/Oz34Ej
yrRhn9WLSy0hj4zHqBQmwDjEiF6TYQf4vnbZtdXvWqdq1n50l0ePMAEe3WhWrrur+D/D1QoJ+RdZ
WrJWYCI4T9z54pc4+GOEBeEJVWvbqQS3xBc1vq1etvOKXU2Lw526AhRTgHA3IenfGVhuHt0D+9ti
H/F1HDnLTJzr8SUjCNrN36Lx0WLTfOsoxZ+0VYxFKkb+tu3oMF7xYuqyvN7TjqqIh31ItIHJSKMI
zuW3VeC6UekK9MKnEY1FBqTrb7CWzPvj8CI5dzzRaUtpOuNQ+AxcKylUmIzP4+JK/0pai6L5n1yI
mZ166+GFBddTm1CgsCkmfGGf9uCz7UXmmqlb7VzklwPkJ5bH4tbGvQVmUMXATsk5T2vMH9gKhqBp
4ZuoAp1Ye76f+A9vFw/nAJDA51wJ8/jDBw7G9mzCt/jh1cxSoKswKunSTul18G0Qlht92ixfWB2Y
Lzjo40oKP2qyJUjA+wBuvwKtwkPobVwuNk89XGNVLnbzocl+XutI9w/vgT9/mbTHLUSLWOdTFhrG
7Ex/V+BxngYeSDq+sBgKK0EhPGyc+NN10BD2q8zVPuYCyeKacp2SMy6m1BR5m3r9W5gAmVOOJQNK
hzgBLFx5SCU8PO3n6wrfjPemawu6SiiwJNAETW9zQWUWTNuYcrvsoqd6qDGDETlT+OzpoKTquZXB
iI2XGrkPjjt+Y1sEbHFl8338iedEvWNaAZA45kEEHZYGv6QS2lv9TD3U5GcpDLdLs5yCmQfQuh8u
ujUD/LWiedsKMQfBgLG6U7U7UgqYP163anE6SgjxwURrPI2rDsJFdMg7mURakjMjuro1pX74nLIH
VzPZZv5iADZeDBbGZUHHr/FtxX+GgM3uJOWag2iqAequBslBGGolfvASsyGwdRalvFkO3Xn2XTst
V5/HQehfsVR3AQ+6hI3Gk3AeU7GnKxOWFUojTr8fBMsjVJ4DlsNWIq93OIZaqHC0nUiuFtT8DP81
oxDLCzu+oZ7hp+h46owouW6FvaWaTthIoZyaJKoGgKU3VuSnNs88LkRuo5meTaU0B2FioN298kEy
KMYo1TmQDiT5gj8gNwoRA+voIhkDQLitzxoNq42m6p2zYbWT9KtHdtLBLiFwDWGHuHQIJgboGyWt
7FAxPgnvoH9XKYaTX3QiInG+zGRaOYFuoA41xpTmM4rxsZrJq9RUIH1wF0EGzxDyw1dFR3R/BbYb
RYHw5ATVOYPMbp3RboXy5R2jm7w1ymIAN8tkMWfpOUGUdbW/pU4WrPy4saZmicatbArEcJYkQS67
feDjYS3203yLdWmJPJLOiX0KrQsyNkRSkU/H114koE1SM9IUxzJuL9gicVilxXWOx5JyBpcUzV9c
aPRPVhCXfoltJCHDhY7HOber/u8b/wpvvsxzBLOYs22eg/TOCBLIrpZBmCIV4xr44Gwxu+r/pR0k
JtY570RhXEn295PKb9Ew1cbjVbeInmwkfMBDIEUKO+XhjTkswSfWWGYJ6F9OXGKKvcPHVTPorZp5
nGN5eCZ3sD7Q3DGduTKi7qQRkqpEiXw7U2olI07aesZopIL0b2Hs0kxpO34bJH/o5jfVbhTGMQhT
o0umRSQkByA0SqDHcD1fXzE8uUOqnBByA756jzfiDHNQUSXc2Itftb9tw4GtKtQCZT2nBvWT8VAa
rtvMmsmnaDsQ9gOJD+NbPuVZnOzb3sdvOuBEvL2rQNZZHyiFtC8SfGp7tM4zYZ5Opcr1vtHG6KMN
cQgyegWd/LCz3tPJsa/Sp5PoIcUai435zRL2dh30FcpISU+qdi6ijA8PZeNGIqcJKdG6oo+tsJKF
rhAaQ0ZYFXe2XDetW95axiZyqSnaNSOv6SFZXLsRPu+v9Cxq/GBxWmPjNenuAZ9YXx5KALNtovLZ
NZgbq7F5U3cQrFYrFoRKhyXODdhmvd166z2hA25Npn+A2cbDfZ+/12TTlAe8nKRLtVFBWVO64Nx/
N+9+ifdw3jzId5it1Wtx+QfpKAWSnJXKTANx4tt3LjMa6r2nwh8BIbeZXRYPdnvEX1H+nPS8dBVO
+eNJNCJeU3CnWgs8UFeQ+urXI9BE6oowpa8PyuuI9ZnbmunAEzdzHSvQJEYI3dd4QK0+0fWxltR+
vMfCXavp2YX/CyHswnEU1hih/dQ7QWAhujLIh5+b5CgEHr+EMgqwWRJPbpDcF4bDEQJHLmzmQZCI
9EHfN+GamyE8A9JAQZDC2pp85ZeUkLjaqAOTc0DJLvzYsxXMPPWot3pvuXZTSU1QKCseNbfQuunr
aRt5AaAJWLvjr465gLp13obodmNxWqMEBDF9oKowx4SXCvz1X26gwVBrA00oCeixWcbVoU6FyfpH
Pf6eIepyIuVs0OeXePtQVT6M7+xaJnkGTTDjdwNYUlMDV/tqzoRvPohcLxA8WdqPZuSPbqr6ifuf
SMoWCRzRfVI2qjkwK5ZKGKTuWfTAdMl3vSn42h5NFXAYDETzW1gTDVT2eXeTuk9DtxSK1+W/ec0M
cxr/pm9JsBkz5HMrAJPTXd/UlQPA3VOvDoD5GIx3YOge6dfLkvclZnr7+VE/fGLHNsb8KFApa/yr
VeDYq8GeRaAJYRL7tCUnLePjoV1yS+jC8xx8AecRRMbM+3X5dajts4mYZ5riJkqbt3MYe+Atsh/Z
KPxJ3MmNjoBCxmQf9H8pz466n3DuFykPGU6zRsvTagsw50GwWe4bAhv6bRC7o7KzLPihRx8OhymA
umCnHe+84pmaE/24eqVW4A26c+O9eWV/IoOVOhkd0WFu6VfmzL2pJ4bO5VM3IHOfiuJxINyI0dDy
cs3IMb9Sr5qMyMrj1H7dQGHHfbYFrnY/leZdH3DbbvCh6EZD+fkyGsY8GFQxBWZNQx6Arj/GheAP
Crmf30dMADQzUyQ5M+znG4nJpsEXF6pEYjNDopABy1QgItqdY7KojZ2Jmz6OJ3emt77E4jHkXOEn
Mxi3yNthvbfeqhDAemVgnlvzb4TXPJaqAIEHTCILee4W41IK3uAjqaeYqFhDrOBgxKJ6EB0P1YzH
M2FytMmQQmNKc40gahSN0nwe0esgvid3C0aP4mZMSwSVA3+VaXOdVR1g28Sv1taYOMfchdrB2d+/
BReQV7nphmFaKSddych4TPeTHvOaDMnc4EuMNLk6Wfs4sgX2h5UPoIZ0EfvV5LXIsp8GQt8thjl7
b7qwpam7oa85by/ij75/dwBplQdYCFtfkQXnanzuAvIhKauonNfURD3AHPet+x0OosowW0fL+55V
KFbISaF8/jKLMny9ZHqTRWo6533baa0LzDMNvDToKUFcG9Gj3jeCXFhQOxyL14um/wM+pvEhzMJa
vU85oDEGMK2qVnZKW/Ae66FTZYkWYNlu3nwud2Y4psqV0XVu6FmjhTmEf42WiXKpGYAbu/3uZb4a
BDavp1HujvGjVCqC7qQT34UhPz04H9Tq34E3EXZjwKhpk8FbxezX4ROB7wuDCOSnvW4Eshowx/cw
UCZdJHdMq6jkpMNI1G9NX81ysh2E1pFIflFNFnYs5l31WYjLpJRjMux1a0dv9geUGNbOMzmc1/Bh
xGH02q+9bZCgODs4ZPf5G+hLJEA1U/0rarXgZRkKOPki/IW1CNQj6bTirNe3biUV2ymMYXYUHeqz
MWIpJdfJg0GlLclOqHl17qQmK0R8Md3eCD4PsS+nMEi0s26Dy+G3EfCdQ/E4XDu19Pf2Qxz4dIdm
VaL9guNNok/dqwJZ1QuLeXRv3wH5aKgalNAyUImTSWcB4LUGw1CNUSK4/XF0SgK6p/OWsqHgzDPy
RGpdNOzqwwclpY+mmshdaa6R3ja2asrWNQ1cYtA0TNfP9T9cWh3WmVhAUOQqxYG7xJxEIdOoIFDx
1kKlOFFF1YiTO8LWyCFfhuIH0NTNMX2uHAftDLpNxlfTvQwfOjrR2sHE0o7jrzT6J6zgfiDFfQe0
ArK4r3K9MbCQCR1xrrBjmVERd9/fmTFnX2tNUZ1XKEaRWR1Rq0OO5oJSov+mdDgfXOU7I01+AsTC
JlLGBo15dOs0Uk8AEdavL0qvU+n362vIS8TzgJi1oHCQZfEawxG3UGYLwTs/YZDpNFOVtq1KP7dZ
GLb2F83AUzXTduHEG8RQIO1rpWLSIjg68/D0pZbbaC2Zk3Y+VE5lMbP+NVr2mo9kAoaJv+meO+cj
wcst99kk0qcx6v/qPusTtiA7cLzn4PVDMflCNXkH/XNnWjsoccHUnGlOqOFrRpnGJdbnMQS8Wef7
Yy4cnLMfnjeVLNyfChKLjsXjPlXeW2AD7XuGbJcepxcUy5sQi4UB8OW8CuA8tGJ/NSe4mRE7Cjhs
C+HwQ4drWAy89SGlpOMLeRI86UEM41SY6impSjVjwpyGzmOWNEiZhIjxDU/dVUVOybenZWhvbncR
TJhC/Cu9dIIlTKZV/tYN/MEv6Rot+QbGFqwzchvQA7KEdu4D3izzWkmR5+3FnPau5yAiei5+hWNq
nqrlGbkpkEFQ9qnlXaAE7GqnpaUASRfBxiqQlv51QcSiSXTqv+zTQ+kSLBfmFpsXX9/GyCwq5gNb
bvPXeIFiSi2c9XQSiltJM/gN3XE28ib8vqF2vl6n4MxrnfzoabFZUFyIOuQHh8wg348fNmDjZX/j
gsV6j076rvh/tP7kIfpmZb+Wa3JFqBAXmptwYaEPtEAYrTwS/e1hIHxd2nJR+KT3mCWIhxd9Zqdf
Lg56cY6qHvwy7v2LxgrkVPjpEPhpLU5BDS+XNg+q8qWdmXrZoHGL6HAKWv/nXp9KGZFJqd5Bx5m5
sNvNacZH14/IDMoOxOKfib8g/5uBfbMQ7NZxtqOfSnTgQpei+AFpI5dR/1fiuR11HO+3npfnvMwv
T8ABqSEurmeSfCsTHH671A/bliHX908R2S0NFXF0c9OyM4birjS73AMg1lZmOY3M35bOd3OX1+eD
QawR4aek+YdCKDY0yq/qhC6jHCf0yuFBuRo044vdsBU5YqQ4dd6/d4P7/3uQj511r/O8XsYJQGi+
tFC5RMGsZFwXZYZc6+dS1/ykrkiab+83pRQdxvnTsIG0dZwjRsXvv9fLfSlHFBgFz44bnDFSOr4b
GYLwd1J2olqmZcLzc0+VDh8NCMMNPBWfsH7xuzX/0rDpGJ03Uxv+of8364kqF3RT4hj2AHh2IEs5
lP2I6dPKfgI4o1wv5+Vjd8J+6pqML9J3lHY/PoSfNAuHz9Kcy1blYPOCuVc4s8oQEQMT9xp93guU
9i1VkJ/+9jzU8cNP9+y9tvUQcFjYR9oRJc78VzjgrTGwVWFIH9aQrxTTTgMFa6BDRW+ZsgOf0x/W
zu9wqzJU1Nuqsz/7EXrwSTKZBeS7SIgLyiBB3Suy5VbOreBbqTooShiSZE+s4b6ZZXmWc8jWOoVo
F5fY7/HOVLxkUSMR1K3w9dyG8a8iq68yvveD/0SjKMg56Cr2K3wopSIaI+uCZi9RL78cvQqU9Z/S
W8xScAiFviZWt9pspLGq3Ls9zoZbjDLUXC6ZkHf9Q6ozEYVNdrXdKWcL4h0SkBIxZl35Ns+er8ir
LnwXQwNn+A9zdw3uDEBS1j6NoIcjO444NVeHk9RmCzmg6TWNb0eFpXmHy/68K2FVbZMfkCPB8cMq
6EuWDZHprXRB/1w8CPO0cAqzWRYbhqFYPuDxTpNm8DdKQZH7YoO0ziKvjZK/9/XR5xTPQR599x9J
yxmTYhWM1HtKD1mSRma8399IEoDtGfFtI3Ts2gpmZ8zuuihChxIJ2QrOZUZiEOAiiLPDe1LhGF/8
O24/s1DNRhP8dh9nUjUxoORf3Os/X0ZVaJMryIE6HqhnyFnkGVKm//dsBEbPazUuGD0IeovRazaw
6L9zaq2rxfpA4fDRSCEcfTju8N0awwPdrWh2YBR1txd4fLm8C6peRrAr6qkJYocJzw610MZT0T6I
8EDI2+VzcuF1PmIwrA73NJPBLdaC10TbOlhBe4nafeZo511HiKi4Qb1yCu98UgPElNAMVSTjaXhC
39XVC8JjdRiPIk3yubhPWtsGXIqE1rm/CDVSkPjlE2BceRDVt7zOlghBBjCbYaFkYJFGHU9N8I3h
ItHXggB4kMYdni4WJwtfTpv9i3eTL9JpACZBAcw4VFM7Pu85nQzaYJ++wfoAC+HPuPpXlMxXC1fu
PzQro2NUxMSj2i6I9Wak9X3Gj31LTUj4+RqXL6xcdmd7EZk5iFhNNUDBL0tnAcmlkeUKyaq63KrF
dkUUTzIamAObgdVLq7Z0IJzDcnOHySIg3afDSVkgrD5SgOfwrHa6O6+bPlyIhZGLgppS+tMR0wxr
cgSWWFWzkUJMQH11ABRAVY8FV1InKiWKwRWxpqnzcn0bpgRIP5IkAdKAAuDixOSxqqThUby3yS1o
xA0mEFdX6qITmctZeZn3NQK03UcJt6bDQ0pWG/dek/qG/lbKAZKVJY8KpS16YEfzM+pxCZ/JQNTB
4E+LBqStqF9IZNaGsee44YNf0M1kxsJstOScdGbugCGQGL36vqOMksO6wLvFf4VWCa/3tz6u3Bh6
7pvoGeGibIZlBr+gugWusK+m7NyEycj6djjozXORGDzBOLFVWtuEFMyf39htyhU1JmMoQeqsTIf5
6QehFvmiV/QEls7i8LqAH44yVDXs9sqtHRD1sCEAYulAGR18Kpe7Nylh7RBVOwnmrGbKPYaAQ5nR
v7Hrlea4H7qgqnb5mAKcVLs29hx6ZszkEJaxKoPc+VlDK+9YFdMTD5HyW7AvH+hjv3GEFV4V5Azj
5Ukc878YvCPTo9RNQRN5XvwxFOBsGyxcfbAGpc8BVOYaPINe3OKsUugcgBOynBH1XXYVw2umaBeP
APHKeG8s2Ds501rAE8DaCfA5VxnrI5DruYiJQsHzy2vJTE8VHalgznEDvignbivO2dR4MmGby+eb
1df2IyJLdvZjpQhHRBdcXJML1CxKdZlX70MNlfzZvmho/wSmqc7yz15NnQVQZqDFdGdSJViU3p+D
PtQzpGRT/Fsr/PRZkMPB/om+ottRqzt9pH3h8WIGrrk/sd1rRB/KzspDh42jBozK0PR7wwN8jZ6D
wGGggm+XXkrYemDREyoGPSvYUQS+VICGppDbWv259Ze0qcYmdU+dd/Ss/t0y9rgnpQF/ZC+KkpEG
nZyYjS7fbggfDA+a/fTdfDB6JiTrC1cmNIHLiRIbAFV9bcMHEcsTR0MVqY+OQB3sECw5brTROL6V
t/tMC8118FVLdQCMuo2lN8o9w+9/XcVdOQO6UoirvEX6/6wamFaD//Bq6Qbyp56OUKLHK+HEMMhO
uPEvI7n3mqAgxu8U8ykIx7brpuYWUIcyKmSgGYb8XxRxjlVTTQ+hl851jjNUUVbN4I4jejYbq+df
FTti2RGwcQdRxlAvE4lZtPb6SLySrp4ScxCg4F/7aTJW0fy0Ok0vzofZULMc7teQNLr5bBc6Rjf/
dznKkj1WSFXv8/+Qr80kDDhvKPq1xP97dxGIr8WsbMZ/ri5ircsAcp7Hhkh6umUBj+XaoCAUPnnx
eEx/1/W52ZWc7b78oQUMLfZdA3wWrnhBT5CgOV5bBSpKpNkQov66DIme35ZqXXAbIZgMl0pfsjzL
c/0BWvV1JxuEa8g6DeJmFQjtmniIQUQUJHDfn5niufxDTrECsEaErIC5NmSqO5l9JAN8BOfFElZg
id2HrxsWpxiNF7Q2kjFjmqsZhaoDvEWWuR4mzjAyCGGlSk584eIkr68fNxYmc+RKADp2++v/0aL6
Cnjy/ELIIqihDPksHoBJd+kTKCXil2NXo4Z7P8gJjrl7VusBcvM589OAHNA85frWY+zLg8zUbCjQ
mMlcYRajPFi6uAtG/UN++qR7nGAoHSB0MaIFoIB3xFQVNNNaiQDGgtTB+wO2EJxVlWG/lwgXfkWQ
vz1IaemnQmiaAE/FzS4yLYRpbsUVOvmb2DPNLLuWkOdZlyxObyyh6MYk8Ql/RnVk6M8ZxY89aTdp
yUT0qRXB7rDsuSSthL3i7Q6bIEmTVhED0eh39tlf2IYhTvBSVQUEb2kFTzxzPzoDwNgji4UaMeUD
67US3o8/hjMc00meTFXtI89g6YMhfVAh2XjllSy2nFH+g/j23o2y0coxmqyVUsKSR7z+gxs9nytF
OYho4wFEIkre2eaHV/qyzP5+jCc3hSt5riHWw/Ei05crGfZmyrOUId5oHBdr6I6QXh4wJWFVB2LG
5h0rzH2XvoS7hBJgzuPDnTACoa3j4glCyFa/ALRBSaFCMcJ3FydJ10UovN+/R9ZHnNsdA9igMB3a
opG0pFV939kbvfJ4KdnxXAeYtJQ+AmxNMyyJUgts+lMLxGGiK3yzZzcPeM9sL4VMM0ZzUTUgm5an
5Hg9xU2hiU8Lm5xFiC/vl1movkp7X5gtaFSZrnA5fEdAJlbnGbHTdriVdiZsV7QqR/GE9I6OPu60
TyUOSP6qdkEUTb6pLz99nCCiUbp1oxBbZhTq72Set44p5E0/nfZ7BUrZ5Np4fdmRcU81HTX0dMw9
yl14y/YACb2IZbxuvnN3jWIxMNkSr1CqsFB8XUWHX5JP/vcxTVF3T8oRw1aeyUoui3Zv35fpTBzQ
w9myYupOczDNYv4UFOD00nI2O1XpVXx1RL9udKN9KRZFDYhZejmSRiC+cODLtvytbi9BKSrrl30i
se1sQF2wmYEqWHW9ytOJwKFISsBWE+B070txkk6GjKJfs6HDDQtSnju+UgVic27sLDw3pkbTs8PN
+x5ispJaHe2e89QUmcxRt/Eb7qxdGnpYK1GxO55dC2EejodeKNOsCZPCC0pKNaw+LXNT+Z/yizXA
LpeiWOKAnMFaxZFW2ZmXuX5uIuqFxNj4QCjRD0jwAsgWL8uxv2lTFTSygW6pr/gZtXmkOwVV6Byp
5D8oDF6yFKa8tIwaUhrjdLE2klDIS85xuLBGWDmU3rE8X1ZWZwPyvnNUW2FJhb96akm4wkT5ILRS
ujoq6WE5kLQ1fNRcNooYpGKSUw0sffyDYk1axSyd2uX3aBeAIRMBV6Ra4Y96zNAToc2mOPfanvE+
nSUEdTMLaU1QHt6e+phkBx2YN0cEed16/LuF1RWd59iBWcJMVYc2ZvvNeArZuFnyZIeJGDJ3W4Q+
SEZ/qGCb0yOS9pMeAlVvvYxNN3I7befrWzq2UDAaMssGYWVI1Sk5GdinUr9vxA4FXH53Fu6VyFYH
ryGicx5QnnhZPiQIJ+/1ghxkQ1v766y6atgEAnQrXLY8FH0qJAjTzzYxBwdaiOVMRVUmiGICFZ+/
TfSuyzLVqbCF4qPWoMbMuCIcYhzQRM1gNB9Lb0Bh+VgNSPBydLHzHzNKVTpriWQmaHw2IwAvkhQL
25Ac4vLm+CRz58JPZ1sYn5l4IgdA2e37jzwvcaKrIw9L2QSQSAUEkw8SBCETeaJWhQiaYr8We+W0
mnf6pDu+vs3/8pq9PVytnC6QuDbLAaGY2dq+h9vLngUR0PZtIZmDUlMtVGFFFIX3LUxkmX54Yb+z
ORriuyyS5MaC6AZM6uUIAkpz8ojvhX1IvpzaNOMuItShS2UOyeeCpNPO3NYIWFVqXSLaR2mHs2bW
+eJCmNLxWmR3UD2bdE6ED+RcepkoCcd6lxDDvxxezNNWkPxCkHubtpMowo4Iz/mCTOvOSIA6YHp/
tfEmUtWVnjpGAvjIUQoVM8PhswojR1yE0NgEEO3PtUlejMsWUU80n9hZl0Df3s5WfP8Sand/c9/1
s6EDv6FshUpgw+7UjIoemwbPhTCtwxg8Pba5tfX7FAYeaHvZDKTNAAAUoZiSctchKtpQ1NvuErLU
1u4K026GvVpHfr6kqznEnZmym1X2UderQhCevq5PgLfloUrwqj/pdxzyU7tnw1J+haTb2PqLnb3C
61dyzECOCo0F95wd8T4C3232n/k+r8miJkREPKVTP46zy6bET2uXWYAN6W12YZXBZ6w7nCZvo4bC
h9+6HMKS3qmMNGa+sCJFmRX/cGKmrRsGnYNhvBtylTzcVBOt+X/bFfYYKwWabxqLPpDbfmWC8LgS
6r/pycLbH4okQXnGKeCR2RbObN0Pm4ALrtqpbo3YiPSczQqyAFbxyJs8t9xXfzE0p0GG/y+Dygd2
JoBQQTxVckMrc4Jmuz8F/4wcu10Hog/cipxaoG7haEeJfXWJJ8nLnMU/1ilqvc/ZlGBJj/wluE/A
EVO1CYN6KlswHU0UK6u08Yx1urdsRCzHhOeEb3cZiGSisjd+S+18Y6DThvg47seAdTkE8emteEyP
OHN5b3u7xyEIyCKnvXZdmEAP3NhDmfrLxy6asagYbjPTAAd+vZxU4H3zoq46G+R6prmlT4PPcUfW
948ir0IZ66tXqZ9HEaxP06bAwXXaSVw3DmWPrwgfgZhF+/1gCwvHDw8E+V0Yn9qKiQGvo24A8DCz
PWWctLqSsKQ4uVRZyQix1kmPEEW5PPryqmfLoxUO1KxinyZsgSbFid381JKg/aSJyNokGsCYbbnM
cqBe4J09BFR2vyio2HIkeijW4t1FMKJXYzbZ2MRirr+ofc93SAjvfG+PpUqeWtHhh9soJHk9inHe
eFxGxLvSWhWvWMtIy/kVfHRKbNC3Bt/M/EK9qQmU/Zz3gSmIsRnQ5vfgeb7kcTeGIhgoJbLUpAYz
lkhfpoFTnAZtXbpIUZygyGhOJ8FYVyp7QPp8pGOeD6BZt7ojBKCiEn9zTvRYppapWUhmg2TrKrNB
uwSip8jKa7A90Tn57Pra1GvwA5jAN/DQ97TnjMmQ1bIAQjwX0KM2ffblRhoE2GcO4hl8VK5PnSlg
iIcPt8f3xN3yDY8OBeiTqhnVtB/x3jQLlmmS9OW5/R6CMTF4Apa1s9p9bI/Jy08lgB1tGwf0n8PE
sgLXK+qPwo5YJ1xX9Mra21TbG9/8z5vOylX5vkCbxp1e0f0AHOTdw06dCrM3nmJMTrSIT4ZdXBlY
PifY3h0LuMZb1Ra1t6CUbcD490N+fbNbXqT+uAsks7SbmW0Gx8HizU3RhDQeX5KLI8EVZPduZLbD
tUWl3Z9YeZDPHLzpebcVUS9wdi88lBiJSTi9cgmtWF9ktN2phA+X9uhTSKgPV6o94GctuUSfOUVU
/8cvOoGEkJhLOrrWQ/vpr/VllzM5HGfrG7xdb9vKmcM7pqMW641zaywA5uFvX29BptzFwjIn+dlb
ZaOk9MCDnCnxuj3oLzQBnCyaRx0IxxqM+YI63n+KKZx6qFMAZJizL7VldtGbeuIu+rV/51OvW/be
stvB3DEE1BFvjsUy1y3RBa3VwjLAp8HCoRZw0SQcAjLjkmd+CNpyiL8tZtaLaV2DIqlRwVJyC1HU
4tbKssdiGJ7tVW8AJKAVaAzCwLyYZoqHN2YoOvIrO81jRLq7W9hM/MxdLoiIzFhHtTBNVwrsuAAP
wxXh/XLRPZgXmDcMOOdoOS+iiNqlP3sVWNF3eCqSrv330TcPhHc9lS/fxQszuNXL4nNfFTlsLVIE
IGZ0/ksuxrriFrRDGYYBJQazMOco3BCsrmxQiiItsJhlU10XyloP+CHkTLsHa44xx+av1+PGmOoW
9OGcaZz4pzj6pTgmrL/6+ZdMfZvXCXnPvfpFiovjASNPIBIW9vuS3eFU6asxMyOn5tiRewmXBsEc
hnUq0pEQNW6yDN1+PAsmcIIpZbqkH9vp4hX3wYND+oe1gASqw9dd3Q8coZBdGpclFwc/8c8bviAy
X4Sj8Gy17uE/WACtLKExBW7IqxWTNLpSt72cRLZa8LpBawAdmeU/wmfhNtyts85wsiq7GjB3l852
DaLI21xliEVEwz6+xDKZNg35NCQK70ArIGqdJb2MMoppXkBYFZx9wa5MCvZ8S+lumR+tSGbECw92
VR79UYbrZgCATcvxJ73PFD5kXBoU4+T/nm+7geYhK8AkVPTPNfoo5ETbtQoAX14jZcJi23t9Rxdq
uotxoj0rWVaBgvghlCoZW6MjbRvPDMnsJ8np3hHFkP2XoRa2QLfn+Wl5knuHUIRdR6OhGL7rei7M
qK5bLJLWgAeyTj3n418OCfGYKjq4c0V95H6zdYYv4zheE6g9mjr4znKFfOKQO3k+cDVAsyUEVWK9
MrDtRisumBdnaUbdO3iJhXkhw6rw0skxdF5IWqX4arlCwxk8xYaMydVeE/22lY9HqXSVAd+Efwa8
2k73EjlkIiLuuZjFU8J2qokAGbEL1O33Ox3oQdY97spUY27NKdYlj3gEU/qnqmjTnNPo75QT2UEx
vJwtFPOJydlBEZhrueMi7AG1w58CVKF/RfHWC1rnLWJcznsLarR6/EQT3iy1pns9RvhmV8CjyJug
zU5jEOeszTfjJmMEXbtyLI6z0BwDRUAdoHzVZKc50XiN7DQ/o9D0EerXj4z40TFJIgaYkKhUyIPZ
oW8S4jggasng4u50k/OTRf1C1wti5KyL9rYdAhO+iFVdu7qPdkZkcwZ7wC6b9F8AdeIfZ1894250
kerHYsFNFdXGd2izCSvMveIC9ZxOyMFry5oYnFhFH9OvkPytbmsVx+PsSAPO+f1VDOPXmK1pDPNm
vLHIVXFjwoSZ35zt/kaPf68nynpPHSqYF27QEU1GqZYCkAPU2U/2EzIHbVRQfnTivG7B6btn5+ss
fliDmzsp3IeDgL7WcJlMrVFDL8COukKrlWHBSNbibm3pUHJmwga0zeTcmU5c2bLjciOYvg9ZE4Fu
e3dxFSn7eGh+EsFYGOW8DceQADFdgRt4zQozkAXmlCHPi0HCotYkMMUHrKaYbPGk76+SBUdGu/ba
gXEpWBlur1xs8dM8hSooxigxuGfxSWPDiN99YqouuMmz803vG2/nEzXF/z8Kqdr6/bfmK1obEzDi
5XNXU8bpipkmd8PaYBJnItWd2/FNBR3VvrQiGRUz5AmOjftmcRVEqi/287rTuylF5EXmwpfWKXlB
ZjMLBwIO/DDY5wMPBTTbMPRlAbS6ywja0Xf8fvfo+Q4J6CkyIZdH1CwBCgEWmwwPOfGPRpGF3dly
qqnsbxuWuJPPmmonNvDGP0G8Q5CSmu/M83JVYft+CIJSdN6s/lW9NrFYaSyGIuOjVB+qBP/mbJqU
bqKjuUND0FUfAtVXl85W/z8A8zE2WiRzcj9JU0ldfq/ImMOOc9F/SIL9+hJwDV+NVKzpxyxciCGF
r/mC5cFicEZyM9e13sP6PL8vHIsatE/quZUTKpmsfhBftBczdhpOvH/J7sTT6CjQTl9q9lMTOy+M
oJnCBIIF6l0kuHcHVnji/81dBTkKkBvBP1PB1lvWBm9NG9gD7j0+h9GorPswSZQairTn28m+WG02
gdXUOLHoD3xBsiHhIKhuPCGTGamUH3/fHOk7TBBOXj3JGnWAYCeZDOq8zxvJuRkXca/PKsZR3frB
gW7RxA+rG2VeLO8xZvRbehRG8TD8AXb+9PnTYuAANMd9qv7EtSTYOZ3N0WFWkhZQmnt9AMpzSILi
ziJT3wF5Npa3MTV/95HC1mVXXVD99S+fwlUwXuA5ItP90OFc7Ns8Xc/eybShSE5Ng0E49YpN6id8
jL1IvYQOOgw0Hz1yku47R8jHMRXrbUIQZJpdTVrrY93jvIR3r3qzehoLCx9K7H1NC7xXhXqajSVe
hgLlbTqtX4LonkSR9J7IRgXTuc4QiL8OvybLAIv3b7P3lWNHG9nld5cXq1almUg+ue8BYKohpoAd
5L/k/XUHqHGFM4BGmyFgWrjmteT1+CqESlGHgb1Xf7esZBjpbiEeb4lAFhzjvTk2QFzkgQNBGvmQ
u52Mhp+UNJIqOe07jqImshk5x8BmPkr7lE4Mt9cHBbnnQrUuqa0qxjHVYAWGGxHVXrkQ0kQoTU4O
hrPR3ImzW/+p7p5rrXIgDTrIkdLPK2L6mgjmI/hTZZ6qSMW4y70XkGMyTCF+sgGbUV9bYEgqYmrt
AcOEFXo3vwt25QOf2f6pMavkwBwRB6DR7uol+DSIEYwu240amtUloE+aL/Db6O5NxHlGiLMRnLtu
uAd3VJWHo76izNf86072vvg1bs4i0rpxx2v+G0kgJ7vlYtMGkYp3xpW+R/O3DIFTVZ3sOTO0FEM5
VtFlog5Lfz7jAK95loCOGT0sENP4/x1Q7Iy7q5JqE4tR2LNT2J6WuC0nmbjFHctNp6DnDfnt98An
oZ3TRvfQd7EMLtq1UZrJkfbEt3tUPOK7ZEfUepP5vEJ7LZnwcFVyOD2QBo5MqiVpNBdLnlzLLh0n
Uvsza89sT1G9U1Frid6jsHpMBcwyRnI7sxUE1aHo94yrC+PkOyHyfPwZt6stJxselvKP2nU2Fx/v
QspFoHsNlP4VyB+xxSLYmifHuvnFBPQw9xgiywqXeTa8EVma1GbVsMBQCO+Nl4qeRP1PZeybdJNs
lZ3iefhnLQ50KAxmkEiy4y5N3ztYV7O+FkeCs1dy4u5vCW5a/ci0Q5humbsqYuHBcrk3ix1sBKrx
xyvP/ZJlkMgUY9nDTiIkIPIemC7Nh0rHSwN3dVhESA8JypHtSmXaDfcV3POsfw/I10NYuR7DhdcV
Oewh2uhHq0QaZw+jn5khif3/IcHsQnNyNcKL8uRQhuTlWruPDZosQmvLSy6c82QtrgWtkj07m7/D
88CQZZn4kmudET3mfUzg7Ma0DgMIQF76iSgGqRX2objv0r2cZaU1L7z8AdTaMQ+AQ3eEU5Z2tp4d
/IYmY2DY+w8kf5NhADO09cUUdJJJFSSjvUMRVEBy6g1Czjzr7eVQjIsj+ym66mzDrFz1teiD1Y8r
by0f3822uMUSHsPuaXOfpizNQGBE0RDoyqL2GWuwjNtoZirVgDa90ZrxHKQKRPYc+EWcmQJl60/K
aqRpD2dIBI4Qrnp0/JHLU/xeFUw7kyPAZLQwn2e0Wvnz0KJiydo26RkRpztjunYTwhPqZY/blQOV
g7GqE3O8kJyCkbVWyOdiiTavyCWHgv0jIYot9K73tcPoDKcIu8p5EQYoSEAsGSe7Z3qUukv5eL5y
cKn8zuzI4DQGRrNvhq0Y9FGasQv8wf7z+QVn2g0Ur+VwKK5+2OP8K5pmx16UVqUaNlZJFbWmPslE
JSW3rHT8Hd2B9fo+ZvwR+OfnWM8bzrMMf2L6j0dr9Wvgf3bh/BfrtmuAVu0OIA0iHAM9f4bF+h8b
knqxWSZAX/7Hl4T1zVtHMwY3y0qhaZCSzxZcU1z50/kNu9ObAWVUgNFEDIxk6gnIofCxOT55CkX4
6kKNAMP/O97dIamXHYZ3UYKEGlwElUr9jkWgG8hCk0gcXKs17FsfiXRXdaMZpwfQRiwXJe1NauNX
s3wOM0pZcrB8wqq8z1c2Bna6tbMc5lJVG35etKdTlgWJqIj0AAoDbK7GdvHhirDlc/gu5ZoGWlqF
e640ayzbNeVGd7N8wY+gJQT68GRhNNtBzCY0SmsLe4WYqEKfKWsyX5oGSOVSLfF7Uf0e6HH/Bk3V
qEU2Ef7q3huzfOX45E8+vu62T4oMalKd/29NsXT3IAO1RkH7JMwDYHsaG1oMcq65jFgpF+omq9Qn
VVDssDkcPUzmRIdYvWBr2o178XvxrcM+W54i9qTENs9/Y+KK+q8/cIq93yZShSBXgnO05r0LZcMv
jCIyrPoP7vWdmyDJoNj4SbTfexQCtq5Vmb02hXvO48E1KQMfUFYwP4hSsxrguJp8d57zIy09CIs7
ll3NhZja2SdYL5tOTwlXj7ddANNM4E496p6heb+MlZp3zr3pQbfr/8tVmpDN/WdthdpV8rfUVoTV
2MrAXtF2h8gO2oEDq6OYngAkt0DSjTFt3y3AHhVeRAKBwYslmDs24eDWskMP5xI3tCfeDmWbjU06
c8EK5zadj1ELstEYOE1EefzNstiFhJnKDUNsbqQHaOoUieHSTK/6WTnrCrstFgalzPpT3SoksMxl
C5lYulXH9sR4YojoyubZJkrphEPxUE6rudnBhSeZWJZyDCbMYp5KJy2mnxCBSWgXbmQrlSwxD9XY
ATZyJTkerUla0jCA/rSZ+CKlKpgrH5HOyGM9pPC1aYLcRH3r168VgtKi0biNgT4SoQ2eLcqzLd/Z
BBOsN0moKrPwPD7tBmp8dlphHWu7A6fK2R9iLjqzChKCVXZvxFsCb69sARgJTRaSwGDE+eOb3NbB
+mCOQD1NAKnTtaFbuWHzXzAcLf1aAuqrXehM3KlKGT3YAhKb/Sd38rDFHXoQLyol++yXaGvi8ePB
pMp3mN9GhH8FVr+IZsdRLU20Dqd2ZyylBoGY+e6vx05PYNgysXm32X8s6yhi433XyWPB7LlIA3gR
CHwt6IXsVqxRrzp4wKLFGgH9KKcIiSLnAq6Py/HeD9OMIUriJjAwb0DmY3NietLnS/+PKRBA7l3a
Ny3b5CY7FDyAuKLlydXlsA7obL17TpSZvVDiuLNwuyNK6ezWSSLYBnoVstaebYOzQpL/5Ao1fuj4
Ik4qiyPGaj7p1yCNpw/XSFbmHFXha3hVvymVzrvmlXvJ9ZfcVJJC5S0cdT4tmDpwPdGOztWHuC4z
MjG98eScuF4UpfYz+v4jg6iLQJiY6tWHIgFHv1xrlrq9tT2eQlERJ03JBgaIYWiIMp2TUrYq1But
qMnZO+2quaN4CNW46YO+WyLVLa9TA07fF1Rx71f0sMKbfY2CKGyMbAPKslcVevnVcDrabmSbpwsf
GHPNCqPENFJwfB4EsIUm9cvSL+xYIMI4I0r0z6GDs0dnAUyKZRMgUgHGpCsfJ93QM56chSkHRSLW
UqABZNfhbTJyn1+UH/NgMeBO9E6MJ9KUJ+6DSifNC0JUsjiIpM/6OJmuy7U/ZpqI2b+xgsdDo6zd
OCYR9pqBu7mjl0vcHexxPYACrys+6hSUPcJVXTz0TOTnjutcB0Wju2NwEq4G7wYIEKs0Ge4EhRJ5
WTjHV7N4A+yIR7xtLGOO8N8HYlURCEAy3SgumrdN6mSASrNjIpFrAeeTiNjd4tMP/lYt6LM4zdEf
mQ03fh22wFATgUluX/gaZmyggyZH8UDQi9M3UyhjBSsLT8MCGmZSAzZTmPeGaHo5XuqEZUGDl1BH
INaxwQF/Pu2Jiuc7z57pY9T0KsyQvEAretIBV5v25yddL+cdr0k7VM1maYfRh4z+sz0AiqdNeIvv
4WlszIwYEcBXNa3dJnRKhiFLcRLRDDiVo9DN2S4ftjqWBlLsrtH5ue5F3FsvRZ1u/CKK2HwkEgv2
wdUplZF7Ye7h1RQ/Nq/4ZPOZjm2IOAXCURWwPHcb+Z7zCgQtoh1cWxkqCaKWf8xU3X/nSu3obOjZ
z9zcKAB5cO8yOpqQ6y3o7UrVwI0gBO+9yc+Cxu6XxGcw2mYBZe3UM0KQvwrovA2lqJVDyesnFDT/
g769FJ3n0lHtzRVpv8ZcZR7twHJ7ugxeLomFG2VEj40wO9lI0MxBH2qAX2my8X2Vr/GS4gXNQRa5
Ek9uI0zi+oC+0k9TDnH0mhQNfbSPNSHlOAiN3Z1mmVnANICKWUO4/XBf+X0S68w2ulf9dOc1uHx2
AO1o1D6BOC87J5GZ6cvsPzpRBRRO/HZIjPK1VPzGfmjYfs2zIY0U2RPMv0j5jhG/TsgZhTum/s7T
KGzLrxSQL/TWpsLXkfzdqo2U/9cvnXnVRHeURyex2nV76HpEw73usdhSvxkrbuyJbgcj0Ak5RYCZ
Os4mEJxOg4+YW8SEk6Prc4zlP7WM9inlq+e82hm6P2pI5BOeEAchimkdIJ5RYrW3ZAiAvEW/gs5K
twSBXj5GzT1ooqwgkoTNnkRM/CrQD+qfFiODGPH+Y4fm3ze+5DfKzSiiNrBBp++HK0wm8Thw1RLP
LT0UUVdQw+OyPsuJ5c+fO78UCN3WNWnHr+ThOjPEpo/rTB4846mpso1hLLBCFN7Q5R9EiA1O9DYG
i4NtEpII2YEW4gJY9TUvFfsPEZwaiS1c2JYI+pOJ+bWaSDOtBO3vihSYEbY5K28ps4clBbdHwCwa
JMvyr1UVoLY1W4vD9MESljc6GxnPmvPjvIgTRwNZI7QovoFqaUNRvjwO5y9axvD8g+xpCFeWGCjw
F/GtTirVM7LCUzet1fY4jjEV13PtZjqeikP/5BiZbow7gyf0YfjiJXkPO1nyPwJ3p/EEV3CjfsVy
eKEhd3nMSk13nKj94cFYMStLa8SbIaVjGKLqRHFdRa+44sYLvM/gTOrL+qWQzRwrWULtswBQRHXm
ivDaNi02D2UlT0ABy1lnH3zZhAEWkqCLqHc2/1/P/MM8arR1x0tRAsU/7Ah/ubnt1onSz+sKGcQW
/vrHmQbQnya4W/5pLlsETlsaUTzh2Wmg0lfh3KmfG1bfccAFe51uGhxjtQ94nYAu1GZM7OBjkxEY
CdapWa4qsfB/RNPhIFvB873T1UCvbhDUdvo7UXbRzEqg0PdNMS0v3v6mOeElp0F+wNr2fgdGEZbI
/sHQwIrW1x2ROMloFiMcXF2ojLPAOHvqQBCEWsmAS8OAS1/+k2mxDm9DvZe20dg61HwpKJJATHsj
ss+ZrOkt1e9lFpsOTr8/vVrdx4zl+dLuQHb/MsxNDmpYO6Pw1lWBp+S5AUUkSJMEauTK/pDfeB2W
3fqHcCZtvme3djW6oQfXjxQr9kSBjd2aB2VPV11B289eetkYq+LCQuevpBF3UVdm7Hu+MkQ+J2pW
CvMczYm/RIcKIhPYI7M48pmI2dbCuoL83/6jAfDdbV+SX7xoPxPLGF0v5vigQqNON3m6eFoE06xJ
Hk6Y2+4Cn6+VhllpuBmzzZz9Jas6eg+536FCIbi0EeF3Y4tcyd8CqpXgEjIl3DycQtwlNYAlMlum
kSF6NzungkXVeEwevRxLSJj3NwUW6nNGi4ygfQcGJF7kvJlfcp5CFG3SO/G8zt3a16f4/vZnDn5m
B8tjmrY1vLNg4vaeFS7X9AvZ9bowfi/+1X4kOxr9pPfVgpRV2Rk+c/BdzztXoqAWIjVjqOapRT3d
hZWjBjh39KqI40MN9GK52e/JkVqUq79Bxh+lxf2h2ZfJ+CKnJMPBjI0TBDZX8GnKzE6/5cU3nxA0
69uS9btcBXEGKKiKEoBibDRdY2u9DnYTDhIZEixOTlTxeF5uR8n3UhX60vWsAQTFPkVWCVcSIVMX
7yH5PI8HqWeHjVyd/HKC0XLe5o6k153IqcWgPZh83JslAg4QaUGYuWwYoCUnIPNDZWBDbx0pHIWc
GUaK7PkZ+DFUGhzakQsHa/hSA39z0zIbYGIfjiKVowgiSJu/BZf0EpFv76Ibqm3orcFNiAAu8T9w
Qn+kGACboQCXvFQfrrxRA3TFNEPl94BZA6U8BxKoQRNNRQvUbi8hEwoFfDYSWlfGp2vjH3Toi5gR
UfYGXE/FZg/DDhxpFMmUNmrc8Qk8bcibcnMYrykkIMKlY2SyLl3yF3PAONQIUae832RQMt32o8HG
XBd8LfdC11AsoOnzOvXZ/1IUzw/Lzw4KbvxekYLPtFaR9yGGEQOVdqeZ650nlPBF0qfy2WneAS4v
LWkbg/0ibHwYpqUaPtyO1mGw7zGvrmVq/zhZpWqd73R32X1oN33H3BnrIZC/xKNCjEyFIpwgAvI+
cEff/JZ/zUOmu6bfru6SZC6XL/Ml83tYLRaCGvMVG/BGleg2cplqS9zKFomAXfTiXEUSF+MkHUQG
dJMfYJxuNaspELLE0Bl/PrYc9d8xNsKqRpGGIAqILbzYwMsl4GsYN3r/w+fhoAP5TUM5Is4b4uzt
FdE8zmQIyn2s8fyof7NV0z/ifzEaUcZeisJTLZMHsi9O8TcvEMqP2QddAXd6PXA9cqVtdKbR0Asf
+0PhcDPzZobwPDKXeL+qhwIzMlutCrQ60mnuvTn7XZNdebnDBw0SIWkG2Hi8SVu+80f8JI2nxEW1
LUUvP+OpsWikCs/hWZnPHauiHiO3Ye1WGrIUjP/vaQR9UhjAS2HhEGw7+mYrbqTpFSLH9oghrKg3
N1kdSEp3l3py+J8wyEw6LphI1EjVziFfq7H/xPYMgFTSJcwG58zIjGJAw8fCndY4dzX9RVdrbgMp
ckwKFcDftwueNpKs2/YJRwt1Izj6RXMLF7fmkwGpdB7nHrejqM9dx6XbKWWQLy2WQFUURFfqzqy/
8Nb6z3XhWy2O1rVmCtLh7rYWJoUjXfTqAfv8Mm68TPChAdb5sOWQK0vFQBMSMrXueQ9WuXwWhS0P
r3iZl+loJsluPsunZIpZv9gZ5r3Y4smdvfh7uk3ZtLADdMnjDlqecPg1mAP8viNV5XHqsebnU+7k
UEU40UHPZtonD6ER6S24oMYz6wJ/hHoXlUzgVNsE07oHHYBYHwtcpwQZdDQCp7U4IKk4DGJp7yeq
7AV6ABZ9sqKm5OKJDCqc+lh6GjtgCgWKylqfC3+IuQqrBQiS20Mc+QZV5TWhpCsVi/v6N0FN9b8F
0kLhFmlZiO9c4au90NFe+mhee1l6lhL+2IVPkEJ7jdQ5bARQFKHuYIeYiNiHXepXYSGnOreccYX1
JK+vs9PcRWO8KTcGmdLBfSqYAKslZSUSsjCtD0eNbHdswj0loPlNsLjBzCD2RHBiuSX1BL1/5fZV
xYG88ME8C179Th9mwagGVf/4lzjTyZ+OAdLtP9o3X0uQDlMZoXLR0437WBvLNKNIzrhdD+NdCwk7
pu4jCQJ3mRYX+SEpfMwLr7UEwBo/QI0u/2YY6X8YwuTMQ7NN8nya154hN9ZPQVtcYJfNzPKs85nx
zUa81MSnXVBd28ErmwaJlCaeL6GtaGu0y6/r71lMaLAompMfHtZV9BDuh+nekfZXblSfBdZoBVjU
Z1AceAqq0qpFZ7rPnz5WKhFxzOrEY8tM1Rhuv9e/sBoWpguxDhIkm13YqYR5DGt129U4UlgKTnt7
xDdxuSSdnp29wtkxG9KEPEe6hr+Fi/J6eJk/oZRtC/jOg8cMITcA+qzGIfLe9sPpp3RCqKbRBqAo
473bdqQmbFDp4jyIY4fOcsNuGPce46jk20EYhuhsfg0srzzI+mvRSiK7+6k3ttJrN364p+dA7/Tj
aOwvkzSdeatRKqsSvWZphFf8231n1mcvvsuRDwk4DCZyJ/AFnCeKDi27ajAlYr/B61ZKH8GIkJ7r
hTW4O5BkJDgaQlv2RVvWod8wAi6FsoKn5onJYNkEZ2+YDFJKynFbnVcGnH2DG9UMr1ucGVj9+MyP
kIlTHHvbkIJCddHK2T+xEwbwt3Zy4OLaCCgPyC563jSdLF/3el2TN6Pp/NTfZ3EUHXDvX7YhmhJ2
afn7huxSd3bGn6fAydGvNTuQNRNjqGDGaXtBGQYolh7lheh8vSrBSFE0ukXoz5fVUchz/AGZ8b8d
7C19dze+Tv6/D0m/XmZ6nOtpW8WeXImL3Ayij1hLyaglqoyLhBHDhtHN84ifPawa6A/ZpMV7w9Wx
mCt85PLAz2gcs76Aiv98iz+imYhWOt699MfMASunqEzZxCGU/jHV064QghxZs2T7ko2s8uhJH3Dc
SjNRm3VMHM2tUKkPFnKySif2pGnEIJf0/yViqgCxy1e7jjgTwhmfkd6dt+ggB6QmOjRmhb7f3s/N
Q5Ad4wq2WdjCHwMo3dhQtPlnYuIqVVP0sm4ldUVV2HHU3Qdu1ehVg3xd/ZuA946WngU60hysKBBI
k2zl8bMT6ZWmtCNBNspSPiA7iAOrP5g8XrrFtpV7Nhqh7NvPFSzcVUQTkIzeMIGKYYYHTPiSKOo2
HQMWyLxD+tyaPrgvRnXAjxXhRdbxuVszUsDpa4qGpjAvJWjSOwM17W09HNJxJ5PpO9X7UcqpUEHN
EyhlBOk2N6Vc6yhbIFc/oyRILFdxMdWr1/4mTUew1QBeSmpG9H1HmyN1SFTiLuNfmeCyYmJOVP92
u6N2gxfKHSy8YB4CYLj8e1GgYAhamAiGa6cW0hf4FKbIXa2zIIzDeNeWzZyzKPTAKKHBnGO+/qR8
C01UIPT2N67hONFmu6Q8thz9XEeOo2AI96JpKdWsSReJZgLZmfHMnFW8S8fd8tSjxyTepwfdripC
SDiHQfct9ZQtfg7obmH06jxigT/gMCjbdT822q0q8M7Z35Tex8iqhQFEGYgaZEj+Wg75ghpHKTDO
COEdc2Iaa5K8sr/Ac/c1JEScK/3in16SSJ5Zh5/RXBFkiDFu10/CEKI5AZcHkx4C++eU26eGXjVd
6qzQw4QbZQJHHNAEi5ogjzaRmUhDGG5/sr1WhjG9GvNMX/RlTvBFY1XH5/+gXGengWmeL4MXJKgC
0kLo+EWK89UAoWhsnpuO+/HyZqQczAZkk+DPXK4AiJbHJTelWLBgmIWmxuTHw05Iob3VlEqJPAhG
Ga66HOukrMh2G8CkGFWhQrk73lw0CA1qib7txaaKmDlwPD8bgxsKkNf09XujOQRKGX4w3mLBe3wR
xY9iMIq1lIVsSs5QRq6hnrcNmfXtm6frissoYaKnC5Os77EH7mPhFGqqrkwxNeUx1AzG9badlOCt
Z7ScZGw9Hr6vQhPse2CZcwMl7703oYgQIPXHtgiaSp+EWRDRM1EeJLioO9OhatmsMaYrzNkKjumX
uYi71SVAk4aaby+zlmC3PjeUo89NKzNHjHEL4jTl7gCIyiFzDkf1Xg1TguMDpXwgT/K63PrtlxQ5
RVYwpeKwRe7ZhiUYDQ1qyZD/Esw2tF7lg3P15YIkF0x/+VSUf3pJhURAYJmL8qQMjbbFc95S+L1z
h96vARMl/j6VS7s2sz/PCR19jvBTb97Xr6eXORKcKL9x/+Utu/NNhLIVib0/q582YTdBlGYI92DX
l5tDovmtvVFiow1SqNNuc4hTdavRgR/MqOA0IVnynBRC2v1Tm4taMXzYeSf1r49LBY930+DtbwWs
o0tS70kTaZ5t/mTPqZ8y5Yk5ZEiktCrBQHNzDhSG5PDVDLg9bzV+HwFtxKwu1m8n3HVxJeUl9XoY
2RuezU3rk/kVrnTZ+A+n0ng47q1C7kos1Fo1G7L5tBPS4rTPJP/f66LUafu5Ej8vxMtF+yxFj3M5
XQ50MpcpNlUNbP+okB9UeJw4zU4/BGh9Y8V5SQh7XWQ7vU+1CbA4CEb82I+e6N6Z3Y3aBn2GzxDh
Z9vfMk2Xx0wqx5OrtifHeTKVmO5elKZxJkEJgb6LbI6QOsrxIkV6mwfpax07643Opkq7UrteQrMY
GsHuvJCnrGHlc0n5HXKk659KLeHqlb8TQZqYV0lNElinRmjvZRE6xzpICCiqrqAUsdb3d1/g8WU9
0SBaT+t570aN7j+p1f2QMy+IvQTc0+Mjh2kqWg3Q7zA3wlNMHwgk6WwEfqqnhEyU2MFN3YBaS/7m
yI4ApD4e79/c91lToe46TOzQ0L7SGluh5Avk6edw3oORWUspYP2mx5ki7Y2KzYhxCglk0aRkDYCV
VyCUWKJjd1YNPWKXcq4mnFkUFQZoKiRENlBojCbtf7m3BpBMTw+zXTjC6YOl3zDKGaGejlxYlwQo
SZai3Ig6Fnt6jqmUdxhQ7VecBZpP/G9QHAR1U2LJ0FSIMHuYpmM6xUi37z6HpsqV8Y8QtXx1X5Lu
Ts7vsFaOm3H4t9BO2xvjMergtEi1I8AHSyUgnQB9W3WGuTlbvwDnDk1EcQJfDpArzoAXoynNYLj3
eCU4PT/Naa6v0w6UHqH1sAwTFz81O+xVXUHRlrXoNSgCkFwPk68ls7+9j6NSUPnMlHSA264L5289
aHMnHGf4q0yssdBKgLB8UyRs85v+Wj+U/x3JPhfpM3mFPEzHtYImH2QZtuJEm0CuSTpm0E/rmyHs
5x/ika/CDz/LEH6fR4q347iQeDlXVvpY2sf8UFUj2NfUTduCkvvaR5ik0xFzyGSjzlF09HgW0g4o
GHVBNeNjLabaEvGayA0xAWkf94ecF+eCuzLFLNBb2hO7P4o1pe/PJsRQ2U1ARstaegHvYSSIfJIb
7w7UB3ZI57Tn+WB18fYlMi3wa+rWwNOUu6sIjuC65VnS2BiMz2b2bLpZ2sHbKCbQPoQd6Ichw6g8
FD6KL48DPnbB2z5IpNpPnhuloV7gImlYO7AdB9UfJbvbKQMWl4tCh/aaNG6TyfNZrP8W4mMlAH+7
iKf7gb/UQgGRiuO8fMCWptqVAettM12eM3ZjhL5iV4Dm5AQx3R2NI8p0aXZwo13QeR0N914RM2xl
GYHKCKH6IAqMw6YuvPu0McLyCY355Q82O/vRpTGBLkaNVVctJ2U8TIDiUHHHQVwIuvWWYFoER0hV
t2Atv9Sepm6BhMqIJedUPB9jI6gYsosW6Q89HcaWzlJWocz8OoY6vd4h8eNgLZ6mTz9DGK6uZftV
veY84nZSoatM0QAiWRIQm6HT89YlZLD0/4oZ/ptAmT5V8ufby4wDhx17MO/U3ZhexuSpGXiYPxHv
Rz9sVqYgDymE4NYELuaTvJ22kVT5msLdptCIu7Bb1UPo94JZNzaEX7UaDI0Uksx1VJgoekYRTQ6X
38YavPlVhmrbxaRyyUnOvOQDR7lefoE1m1m5G+IG3a+rXpwxO/OP88Q7PL3Z30m0pe0m1X1R7qs8
JgAzmn3244tedHTEOuQ3+RFuW5aWV/CUqlXEXxo+0W7yLr3+D4G4Oe4x4AvCgbpjAmBQZKBR2H4X
w06oatw4BPrzHZOuzo8nKTal64sPMgaDyl/dqg66vkFZqf04qFLg+qkUZPWH2l+IBi4TNk4h54Y7
QyrFhfqBAaVFpqYkw+CC/BhTHkRXWQazku6wqm/biwvNHFjDsJOMV37giGyaHp/nbcFMu6K8q7qG
okr8DnFM/d1GRhCtcMBTiTO2/1ozWBhbDOKd2BrzPVQ0Ca0+AQBn3prlTig8KgJ6HhWX7zf5IyMJ
VTmsysHlyN4SliOcS76NxlTmyyu/8BesCORDqM5PYPySi/PCshJwy4EJVxNBFjl8s4z7EK/8U/PP
3LnJl+Ow4H+LDr67Yvszm5rfIoI4AVtVMWkh/AStjsuRnWUNTpxM0eoIgH3P4rvLiqKudUBM6Ktp
gzY8B92hbAcvKeZ2lBSWXPGVXq0AK33xo0DD30fzSRHLCmPgRT8+0XRAlOrj4Sc5FyW06HdUZPHt
oFSZ4/Gv49jwjasmMyiBXWxQ1VpLM8lSI0XP7NagTIegZtHXPHfA9TTLCUkpgDXu+GgkzNzjMPFZ
19H7l9aP/kE47r+TKDioLnUQrF45xVjDWQs5mmh9Sf9t1yqjehu6cZwxB/iJCrpsrgoNwQ5VqAuL
ubJ3Rd9IhmnNXYb7EQSrcWcKRLJK+jCQZ+wNGwM6tEAphQSi8zsxHOWGBDqKxESlJFEU7im76Nuc
BtpyryNqoL7jSFappNA82UJcrTAsSb5bFbXt+GXuEuplDm32OmC5Clg63GczZoMGLYlYuy2hA9Uq
UrGRP1cMuUyYcvbAbhbzuX62fR2bNxO73pCf9OVOEIuLZz0QKNilP68ZKbrbR19291wbATSLs9kk
VZgzs9LzPbVjZE99m/vqGOgzV759vDFEgYY+l5DDNq0xklhEcyFHpMEs3V8mY1kZXZAqcS/HjmgL
94hyHM2iEBHydBhSWz70wuV3VYqW43XSiunPWFfmA2DCl07E+42ppQFHiAJTrkj02v6GoeEmAB+1
/HBBgrQ+s5G7enL+ThW1QkoohsTZK01/DlST8sf65XqT18BIOzA8sCcYibRq//e0A6W9Q+3lfMS5
3kFJQLYMkpW/PvEzynnzVm9qgdYMmJ3osB5PEnJ9fBG+3t36wz3OXE+eNv8UDiH1pD2RjsvKY+ht
sz+tccJancqMuwVGYSkupz9wCy43C/1vcpW3yrNF08PcBOhAIN5tItrgQ9/Ah9wCWTQVaPu/58s3
BXpBo3L5IiN9Hx9S3QbYcXq1ml23OETDwB30HH26v5sjvt/Y7KLlAu2PldAunr0vF7JQbn803Jvh
afpjj27E6RvaXaitRV1BwSXjib1qt+1iMH2JRcjzT4XVUKiEhwS60LUVur5vxmNuqv5z+ISQLJYI
8XZoW3GO1/d0EMX9HfcFo8gvhcq/0mQpfJbshdhJoH4Gf40sMecHmwXVvwdKCwe6dVf6XOfQ3EPu
ePU7/rYNuDUNlJ5P4riZFSvfv1kZVFSGGIGmbUUBwl8JXrxKTGyl6Ezz+/25tGiMSF+DF5JCSpiF
OmMzAGxzq02PR6RoqSIcJbCJBnwyvA71lHZ0EmbtIqdmL8zuLqG/Y53jveWi5o8zpboJXYyqzNgj
Yazzc3eIM23lea+roWMYCS3SCd/i56e4807LNqIFek0vB2MoKJb+jSFyZ6OHT0damYEFDs+eVLr7
SpsVXafgNU7QXeAVgJqMK0WeK9etkKCbYCOpogAOQ8ddSXhEV7ICMyFeUUQkF+OgjVyBMkE2hkYZ
mq2APRYj4Rw/3UJ+TSc+xlifBtzSzF8HOAowjj5KsU8M7KoyQvDDp6oS3PxFyh8ogPp4/2fnv4sh
dNdIyqCYHeTgifKjRvvv3XbWViOPdOafnut+O8z3gVF3KjOnaGD04W1sZhdiGL+RxWsCrZZNcLjX
w6F4JWhMQOXMpcCx9gMT2QtM1g7Lh71UFJm8O6VLv2W+2UZdfYsv3H+c4mbHf2F+UUECt8D0yjG/
aeN6I4EmYjUZobwfBlX14HQVxlmVK7zXrEL3mzZ1O+7foo7QlaP4YZUywVLDxOxO6OjeQ0A/rxdL
FSkAhQXT0jR8iCcRQiT8Jm6+ptnWAHS6Y8yX67w7fzllsGXaD/tyV8PlKuKww6e2CBGggEfh4hAJ
cPNnW5t3uhXgXAPez2O85yit7X3ZxCkWfnWb4Kiio8yyHyyK1buI31SvXByAj2H4YdxNKMeHs4Q7
GOr/EcDLnkiDY5H4P3xyKfVRPF+tYNso0NFrYxPW8m2Cg9cYP8uF3OPzFIfUcx/EvcxU8cLVzCU0
Uvv9q5UDhoSRI8UsNqfEOBDMshjffJ6mwFqcMSXHkzlnX66XurjvCGKDYxJHv+kLliXarNVT+gw0
b4XxbYrsb2/guDpppOJZ37ZX57qpE80w3GIqmSjrQTh+ktWDVn3lHIDsJBYZn9bsiGLeihpEKE8Z
unkd7aoDyTB9tgOcxuyHiffqmO05W1VQjmVhci0bDvq4j5jQS7FxGx4JU9mK/2T1x3GccUtzNKjd
HS/lHkaoxTa9matv1jdrFIaK7+IAEFzRfJitaUrgT5BauNFZ3NKTurwby37ksawJaqqY547oekSM
Hh8tD9Mp6KYpTk6c4m1CsgCN1U2swqdaYdFzUpBlDBi2Aex1HMUIyxOvfxCQNhUUPI5lyWjM5qeL
blpsFmSgi4Q2s0ct/hZqueCEFlhOUW4sVAEqMrO0/EJvJ7WszMsgeB7oiWQChGHfdXp2vIfRRCIZ
MiUYniuYTE96UAIACjYeoJfTd+uoB8VwmilLcobPm439Xbd/FsJzzNvOsSTxEnucAa5VB5K57PeD
k0++7RRJEnDZr5GeiAIf2z/MI8D0mi48fjVQSqrcNxJootNCJYP+i5asOCwmyHFQe3QQaKPqIrNC
VBQz0RrKOQx/y1kfdiQxnI+piWWQ7gtGFolQMudU3lK5GmWT6DidYzVSUYCZmwm/dW4TJHtlPn0G
Gr///+KcVMWjfeNoV4Lp9la6rk35PCCysHFyuK20qIA+wtEJoFAINS+HvwWcNdEUbAO0gwEVypQh
zuJ89IzDvWmfon2S0bA/e2PpOwNrCoAP13gQF5bUNeM3RXblMn+vAI9FAXiAR7E+ENbiee4HtVgf
06UOfMmWOc7WsN3FLElS1I/MkAyl1c1jk6IgYcu/u71xsRGElvPEzVXFSFBhfwgcJ+d+B8fZmPcg
DVmXShOBwVsNSkSaisQ+AwYmQXqPPdEDp77Wx+3z5Qig7jr5cYpsCNy0spuuiND6GNSOi/jS+znF
adayasHl9buwvB5HZFwCElxqn3V9lBwQbfYALB0W9p1lfW7AHRgfyoInm7ldTfBAn5fdNk+68UJU
FACFOEFAz5Ga4FKK4TALr8lnUy1U/Wm1/wCW0sBq+8A4zYykhCWlzfpQ3JvzlbJdZ9JglbmYzLGT
Nporqw7M84999xFuZiuDeiIH7cqQ7OlddVwgOb4KIP2IdkEOqS09gabeym9c/UaJTSD9ypEMG0PK
P13XFhw1noZz6g60uguweKBP7YPQ5Karwp3MuSzPQv0j0j9lhtYdlNULMOO0POTv6z9bX/j9X/YY
j3fjV+2UQNmVhA7pcqYDYnSGpiPD2z+d2FhxDRusrQtrFryaKSKBLKRkOmnMKHChl9AAqJ/gL0qQ
xd9p1ASnpk78NnDLe38j8eAi5lcPTRLYu4LIXzD2GyYKK5FC3+hHqq8c+9wotFKxJHLLVxviZfkm
og2CG+a/p3vZy1m1BYZYJpSFfO7UISXAj4Kj1tMShAVHjeLgb96Fse81f63Qu9+zfvSkXkTUiHd9
nOfcFic8GuO5DY+EgxoaKL/fJRm76iBnsUvnB7x8A7ZyzqzqhLC9wyTde5QhPC8PJjqN33ZfQ0MH
MRYt4Y7G5HVaLZbLEixPIeJ8VIuHDT8d1q1fRf/QWqPMmoV6gLH2vmDsn4CxDVDfeTx1i41omuL3
FJTv0JKrnNkjTqywO0cyuOTyWYIwEGR2Cw7OVsceAxQzafpN27gZIRuOdN0zEjvuSt1glL8E4pJ8
vmdSaFSgQDDl9+d+p16xZ79CK+/Wv8+YR7a+NBLckzae9ucA7daLkzsVrjfuSWurd8d0LTQyPti+
WVpLNAvTD3f0Q34SJlzsis1FFZHXtXk7Hm4BHmyGBV9pIy78TeDekTalwphm/62JEiFVKDfFX636
wbr1Jj5pq49dT6rm9PdugfkLWeViXH9An/+RsegrsJ3a6MKyF78g2EcDh6/vJe1VaTIE96xs0KM9
Y5CfyPxGn22bLNZqsNE56gNBQKM0Xt+tTJQYa3raQWhUifOU4vxsWBpKdCQ8SznINAj4dASiOTMK
WO18XfcKqi5P7ripRm3+niKm7RZyGrLDqTaJzfPJERvqLpV1OpW5ebuS0dUtjpA6o9AHUuIZun3P
kU1tzh0k23PACr4/CVF6g/T6vpTpwe/QHgODDQUTjifxm2XKCrapPmyV4A82keIfn8+0uqYxkOIf
FvOusNYYfvtHSwCiP8rCoF2iaj7zhim+TH0/kmbtqaVCF604J64tQtSSSOFVVzkuRCHBQkYpccFC
BcvwOqGhLISY2J8lKMCOnRd+C6GRSVgm15lY8Uu9dG310wkdpGkiR1PlcRtG7fLMYX+UGyWW07ti
3O+PmXbkiDIPZDcYgkH9cLULlAGdZU75fgqn6Kp+UQb1DTRRlljQTOLJBkSJL4VfWARwHeL5JrKI
FpGeNo9I6FOmcpglB+lk+mb4/ajpOlvsJAJ0TO+jxvKzZf/rpFoV8NaJT/eJgTznFSdm1tK9MIXl
yM8rO1cgg/vKVcvRFbKrPAr+K5BG5UWM+y6HPa7PjCeXy4BMjSA8iYgUKMNuua53ntNXNq4/v0eT
vcBhQe2YyP+edTANC94XVcWlRb/+EsJ0wrnUtKGmTR3M2nbtHLiXBonggn+rKGuX8PR+ypP7nckM
r3f2LLTqZWRsH99anC5toddAj3jb+KEEOirJ3Mgamsdnl6vPI4i2Ddj5rb49xLVh7bd1dpl0FbLz
zrm6kni02oYCCRtddAk5oUKj+ibwmSPIaM9g4pD6vy3gJgwbb0i86sPgbaSyOWtID5fbeSk422SA
+Fcd4f0gxUG4qKTUDtjJDKtwcthl08YgY7CWqyr9F/V+P0YSlyKymhgBz/xvNDRpQ887xtvissea
Dp48htas7GBckOTCf9Qf0slV8Qyyb4LzzWRnkIKoyVcdjdyncSjqhPzDbzkV8pNDYynzmf1vH8Xv
weCUcCRKbCLAFTz8ZpeVHPRWA3jM9xaXeaJEr7rhcCBGc39nUrzArhZAryArERG+X9KDIJ/NJ/0r
hdEuwJuA8Nck66pCru4KwL0L9urP3MK+2H9atLXQWcZ0wpms3Qa/flMU0cE5wJNtWZmmCz3JtMNn
PJkX9wu4h+93BZ32WUR5SVK5Y6HEjnCCvignAKPWH4C2VgsXXj+kpObver+Ng98CiQp9eC6sFThN
F52UcZJnbQg7bax+TJ+DokAIFe0yCdTehfSwWTWSNI6ckHBW1r7XAt/TGGC7u/lMlwtJS0QlLj1O
9irJnk5KpadoNUKNtZ6Lq/PgrIG4Lv8n+ngZkICzdYCHJYYGkHDz8fw8cEB6pGAhq/a5pTRBZn9P
ckimBrCwnvCw4EtdWbpOKXnPrHC4H10C4nkSufBJtse8hIgHibRUL1Z6cfldChu1JOhXUGJ8Ybav
ZqKXgJwcrQgP/9tytPIMqHotX7pDFyRut/YfmI988uW29EZrsxdM+i4nztczxSmj8bdhT+hBNzvI
w/3JMRZ4nqac3gCGCwrOeFhcqracP851e/vWrRYDscZ1ymZPedjPa24mYBd3nSMTQIxRjQDk4L6v
Ad36pBhy22xNLac2rbBKtbovaTQqSi4TLXli2kIWfzi+H6Kr00/B2yKAENiyO/OVB7ymukc4nb5K
ChdXPmIclEXFi73QwdBiLuEPsBUSm/PMqaVDeB9JE6kwypB/bNFKHFYL5UL7DgxlSN02ODpfkdFN
8jfxRN6LeNnYRdQnbi2br/Nmjed/h6zLoVWv7BjQGw8aSwJasHGKsNRN0UMb6ptjiNt7RXfUJZeN
QDi0AWPEvRr5h1LcAbIh5NXhpc06cc5wU0pGE/uSTqVlbBXF5mANKXRJl2ohza/F2P3DeKfW7WKf
S+uvhaabhfhGPl6EruqbqVlTwDcnc6jCEweGtufMu8qQoRq2Ereb/emtvoyxp9sfe+EFdXNMqYeU
tcnm29YK5+/A7aeC7HOKs2Axx5QD/WANf0ujgY4jH18rlwcJrmzMTfTqSG5k0D5eBZ2IfUGvuZhJ
xrcZcgMQnBFrI5NIq/anvIAz8HLp7ZekKw46qpCaOVQIhNhHLZVHEEBdz3+1dvyKgQvihDX22RcZ
mKXd5jpt7Ym03e85USEcj1F3c3mE2oIpr9z1Cl/EbF58AQyJaQ6xbXajLl9jR7MGfX4KHqOat8bw
ErFCKwTcgAkYdhiudc8ZaOdFp95OlYVP0zZr4498/ubwVv6VdUhLu+/6Yo1eRRq8MbmsadVY+741
Dss0DPUC6f5vOdAY1IfPdVq8Ta7lGSiDlbT1u8CLFxHWP9J6F0JbEZo1yXs1Ivxy8ufkDMRNGJI0
M6JSAgyIap8HSHP0HeD+0Mk/iUPv6hpmsIwoY2kkpguJROIp0uSAxnouwE/sAAnjpGqwJ3zX7zju
WS8yQ3pL8XRHRV0n1l4DTTk+0WyH66oSkHGupigfOkGj2W3dpL3GY3URr/x3DaN9P3v/gGFziSAB
Nyv3hRbwiuXHD9Jc33+d69mDp6oCo0u5DfecrAytpznHEiAo2zVN61nAmrWXKDpYTD0hMVYBTvyY
E1bJGQpVEtJLXN42BTOYB2BrgXWT20aEGcjNrDd/MeutodS5C+hiRDfjeU9CQyiBgbr0rYvVcZ8v
knM3QoVDmovpkAXWotsORKUBJdL0UxfTdUS3S1Yluap+eUYIv2Nf2g7L4GQubSxOJU8isvYUPz9l
bRzLWr+Ll/yUJgjpAUz0QqI0IdKxL/nFMfcIj8utrPGYZrWOMV4EfnH5rzrbSQxB26DOhnukCI2J
4SEJa3vXa8Py3XSiTIM7m2Zi8zaCuhfC45F+nx4NiNhCpOQkUJEjMa7oblSlZ+k28J/GDdleKB0b
HX3RgFOWAr5K4MGF83uVFex5OHvErcHqF85m9kNwoNvtNbcCtB4F3MXCe44kjyqG59Vn4DZMmk52
OHiZ+8wtUUnwMJIDHWy5t0FshPUC75j1hp5ENFStzi8mzgUuJwWoTDrn3vfXJ9xep4yTRzXauO3C
PiYwOR55wr1ThyC+FpS4rYtR7dOt/q51Ha3DggN2Z1bMQkx52nSBM7NOoshNV8sz7NAf1H38q5q/
NNPgt6HhHb9bDhbUa3TW/f54p42ahkR5G0chD9XqOTgxxYJoCUV94w4KIH0ciXkWETNciGhSvWzG
cNPdqRxOVIQ7ZeoWlLLLzNDjPwshov3aPRDyUEtvYP2VT31/A/r1f5hNtffpJL2zwKSLf8ZiNENp
2Omo2fEWVJOQP1nrBTBcLSlLQVh6UYZkeAQ0V/X7muS+DRPIw+h0FwzfG22gkF1NDkw2fycIcyUl
K/gDw5ZlNouA6D+96efp3wiuDvcB8CVrI0XqpTnf89KISWtKldvcBJBzwDlsHG8uLZBMTCPtr42g
dgMgsN2E+2ImWN0dJv+Y0tzmF84nxl4MXXEjERjlSLRN3aSBu7iNbF+HJLchns2wzv8eoqNWKvQ7
aZruanksjdkm79ArSzQvyKEkj8WNOS96a8zC9fOs+d7i9fAzl/vopXcFdYoL1dQn7waqqRCkgVAS
U6AK2JQui5HWniI5038/1X96xagRP3D0LAAw3VcovP6fJ4oMev9mTu88euAbCS2knM6A7GKvfMEz
IvUi+5T1lGeqU1RjsKn38I2hhW2tOe2nxcN/66FshYunot1FLEvNlPOsuSM2wZZy2qF1Yl04A3Hf
mC6bLq/HebxO1eljjQRnVJSuZK5A7FBPms0olGl98s6X7efYgCM9v9m2Mk5t+AnkR6RSxsYo25CC
K4EIc97K4sf54MKSGgePzAg+xTVTKcR6x1kssixVjirTjr4X+D5JWTewxsIlJNrk+JljxLqat2MB
52/mKNuL13fpSTl/rAIXzQHaNTKW2WFzcGYKdtpcwFP3qO6G+fGY7CCpzsoDztPzN5+AS8OX+Sf7
eQJdO6riZ8ovmU1q+vK3JOgG9gQj4VPkjq9mapAjaY2kP8M9e7ghyQx5/AwWzf9JsVx74NH0aUqp
WbFZ9CmoSx6JDRkqq1bhp2GEqoRVKPEozXI6lXz67dsbtyfS4ve6rr22YUzhZS+q5dVq95sY2wyr
6ZHhVoRPF6rl3K6QJArdOms3VYpziotOQc9W5sOEqihfb3wSGw7Oh6k5d+keK1lidvJhdvsFzhjA
/tn+jOBefijFBbNMunRWGWGU/lEdDRfen5BtNN1qkbWyi8g9X9B03ejmtRtOhZhzXIdM5Yd+QeR5
0Lh0plH3lXwGEUnNL7+ju7t1j4hpQcU7ZAg2vsXAEKpT16ZhOuCfFgyW9kj7Z9q8lIRysDJE5tEC
QEVQAUQnl4RaZ0Y6iICwjXrg0IRe7TlO2p/TZu4Dmtff1/BmscGDGW/qyWPDayf7LIt905WpRp2g
wS+ofBM794puNWiSoKAnFO3aMJkp7Dp9cYuzZ87tVxOyqDGgGFMp9gPaRavRZGlVM3ObuVvGOWPf
9kxnmYnINvKf1Q9KIenJaFSOFpSHxc5iPNWLqDfcuZn3C/pdMC0MKLgr8MXzNcoUlDkJrOf4M0s9
GcVNdO/e7z+x2/W44Mt4jRRRzk/p/Cxn9GF7recWg1h2fqKYakn4yNtVYkzujIYeFVA1z14GoGWu
g/ndVsZnGlDG6Fr7tDFdiwhqq/DQVQLQxqUv//uZzN5vXHkpxmzRq8YR5SqwCjaJ5T1C0oIHKMnD
7hdXcq5vY7ZAICzsWUfnvp81eyNzTKxiOlx4paa9w3xLq+eVvdoct1NjOGXOdtAWNJn23s/EYc51
QTkH/CkAhGvu1rvGQeTNb6bKhcbFBp6SRVolbYqhtmGsSJtK66r+BnQ7EYwMSqrZAUlq8ns6X2kH
jtFMjVc4uYW9uU76CI/qmBU/nweKr+5/SwOftrh2SufhFKi3qB6VxAW8/j2oezCKrPN1cyHVJvj6
27aE7G6XIpsMX1kkQ5JbGPbbPqZKecLg1lzaF9IsuirtfN77gMSIplpCfAfFQ5Ovh6fLCFNvN9mO
Bab/EZjTnzIKL6QVWf3hayHYEUv1HlICgIbP3FiHExvLNzzLL44kpRCRxLQRYgoIlKP1xLt2VuM+
sKxtblOiRaOhtIRw0eROd1oMvC3WWA6oF38ZZWi5EsXMS942EGu431mtp0piMdEjlka0zGdnYXVo
oFls8vBQ6J6tLKygW+qW85LYgYMo3a1sDPbrXI4E5aJIfFsvehOxoNBZh78pzdBaWDscZuA0PVQF
Q5thbS4dx7s8bAf1CUdIgwykN1n/MuUuhdTptjbUKs69rwivoWNj16N+WYn750xtYE1Sg8yEFTmw
/qkSdHreeGi+RXyr8s2dWMSJ8SwtyTSVUslIwxS6J7Vm5i/NV72czbVGcQTQzniZs8VguYmcNT9/
Qn+t+MuDyogTYDdBk4ipYVzUmsqyvPHVIWc078V72Kq00Wflsqbrd+SyI8oEOsMMlNsQEvp2KtjQ
pqOT/7f+TjuD3XsVcGL50gInZqq/I+IKBEMhxUrRPtvbVYfIx9/YYMr9eLETqNwTeG8p5YHcIoyd
nDDKHuqQelm+RMEZ7uyb8f4EGyoWU68EOHJVpXhAJPurANerKfU8XtDKuUO1uLlyzXxtcx5pR93j
xCQ/ywScdkSMlJt5tLIUEtk7TOlzCPuof8/Y4+vNG5xrhCd51t/15KXgJjjk/dp5JrxmMwLvuiUv
r8yneIoMx1AVkWwZ9AOjQS+pRE5lI0hI7jlaKHg2dQ+RlfFT09y+37KxV7wSxaVzsssZ4cZiy8F3
qjVlsZ1LJ110itEfqtpkodIcc3KynYTcijK0ocmyGt5+RyWPBngdEFbYzNuDRY9HpDK5nr8K1ImR
e54iMw4uRUrjRMaK/V9gw3wDPCQ2CwXqcC9OfUyol1VrpY6CR4LWXPxjfmjApBDBbAsmMenX00/Q
XVm1oIozaBk1WvriTb9pnzMrLkGPBz68z7CX6g8LlCggrMcfynlO9jJjScUGuEmkZtHXLwRYp3qg
dCTwRSY+fm17lH9JoXQ9A7ovXoEIytPJRHN4AVt6d+590bHYwEglCIZ/pUbG3i501zxB3mKsFrn1
zhnQvY+Hj56l1b0NwTZBYJzTMVWXgeTg1LM/xtNtwsoLTk3gZbSr5rtt5InUDhciLL/zC+CZ1GqK
HnNNSKShSXBWHbldSdLoSdw3am3hKQynd3DnTb49LgLVFoUDM/VVem2EweVpIE2AaxX6Tv+/Bb6z
z8yBnKDjhF4NU3ud1Ho+6tE/nZa1HQWxTcy7HDqwnzEttlI7I+Itjxhz+kx7QQcJHgqIN7FSAUst
t+6zEE/gKQ1ysIMkZC40eybucT1aEoRuJNrVVE0NwuwuEyK8/D5qAEba2K+Pc/6x4k9kCq69KqjP
K5NYiGRTyCShoySsxbRdPzLXNO3Wh/YZ3hOtGYdApQY8smujbXmXKsE53kHnCjpR7AtiVdazgt+I
co9wIL7ccQKC3x8hipW9OUkiNzzlOH0yZzAUpmn0bsEwQno1qwagO+XzBuH86SMXffYhuxfw34j4
TC1eX+XPvndw1SV89LvFcfWoXag33yFW8RUZgsjcMs4ffiKmd/a8RHhIH4nDZrYfAmg1zbKojtDd
AUYqMcYpaDpfnLRUsy0bvko3byxuaOhITTp4ianateTO7CHe7jpvqdnFDRaFFMJ3GDR3Cc0pfsK3
KSf9JTjMLYSGL8QiDrRkXlef5AplMIjgXtEXLbihxQplw9gZvlJxIN8NhcjNlyzX651iQUanBIjr
QAG1i4epeQKh4i7zHDbgu8ov1xk/7SjdkVdrTj+yH3V/SefOBC/RPvntTEk4N7NMLZZ52zN2eH2Q
2W1I+MElvkKMjRTO5PzMsOpDbPNvcQoCEz8KpVNZ69W1UuCu1t//fHB4z8KCB8/bqqI/T9pHNEzI
wAu30/j7gZjYJByWSL7heJfTe9BwE02OWqzSZp4BoMheRdxyvc1rrc8zCULRUiZ1kk64ntrMECNa
hkkE9j0bGCjLsHwT+5GAP3v9KYTfyC4CDYWHAriCX/7DhhZEQnsC71jryF9TXsRT9Vvqo7VmevOF
R+MG+Z8JGiYywMdytOFg/aTd2hwem7tIda8BFJIJif2q4KfTAoAslqNjbGLD+evQhbkKi/MCYl26
5HqGBnf7hEYCtRsi/88NrGBdDF+4+UWe72FnuFgNkck71zxLoHSv2BVMap1EqmwQiOxLyH5+fEod
wWdD9jXFi3mkWG1gECmkqbHQEUnehYMPjRu0XoCjDp8DCHfS0rIx5h+zjs3qn7ItyRc6uI1Rnakj
FnPPXz1Nbbsl/qSPfq8HBNa82Ddme3rnWvUgJRlZ9GvuRFLKn5tooFmjgKY2ekUY+ByW4+EcJY6f
p0uOqAGRnyxpjlJH6G7HzACvDyJut4WWFozxYKFjgGhvpI26S/3shsa3W+yH+2CaUW+bWvynqyIU
SgJtnTSTfNwsHK7rUoG/TlELRlbH6RhaLilJGWBQMbIIjhW8SSLakL4HjPT3YDVHuiKMGqueuoPA
pZRa7nvIXFPQeywGxQ+BtTpkexVCV7bsyUckaRSq1hftBOXIXbjQR7NZF4PdC75Ej4T7ssfj4/iX
ju0NKKYuYTLYP/pClqVOUrygvcfjSUhcsE2ECEeoAz/NhhDhG8mz8rKZDD1KB9HnuWH//UnO+n/v
A7l8Go/UFAWs5Ab0WwYYB8t+I7CIvmJUQCyqb/DlvN1a/pqgb+QUA2XDTPWH057D7ZuUEZrObjWy
+RhmIaowqpyc5Txl/jcls4HPhiSgMKU0CNEj66sswPrXzRpZ2kXtn44dQdQU7UoiMWPeIQpSbjMa
86NARDmUBceaq6RT5nobenrvAzanhlhJZu4aTYCbKD0xmNz/ub0n8D3SyJQA0PkwRijiufO9XSS0
8n2mhPxA//gGerX4psLtveYkoynPm81rATGAfWGkQh0c62D5OMh8vbtLVOMlGNh/TigJW44ULogT
VCwW5il60XJvnbV6kLrdXt8glpy4HdHOWBtlEqutxelzlxYiJTok5MerjtpvncUzxOhuymBuJuwS
2Vfj0fLLN2oLlqKDOhbo0BitAb33lQo+Frr2PWRCbGqR4Hs4DlKaHgj+dmyO9zi0Kcy2Uwvv3tSS
9tm/O4wqBKHb958B+50l742f9LLziNYoHam3S2X9yBBeB63hUsXgzzwh/A4/mOfsBDB91Az8NVaP
QRUA4IUqz5Vt8KmToq0HMGHFfS7OJQ48s8+MZ0gldKSb5JobKJHOL3OgU5vW1YzmeYMjgIhOQGPi
53DUaAlNd5JWqj5JumZZ5Gk4zspQe0mkh5DMZOwiMqt2VYDaAK1PLTMisHLQM46k0F3LYSWvKNBD
ChfZSjHmdoja/E7nlxiMOeWr785RRScr9YO+Q+AsA37GgXn3ZTrtk/Km/6G1KBvUIFPJctcWn/Rt
DNSFwPzUBrIk8S3fmWtkMRkxGq/X8pckZUrvhIpfzghWsei3rDpTRhAsHyKbjAH4iej4/sOcqOeK
2xlpBc8Tcqro+JbxLihUQIgCN6gOCCwTwalH+urm+ZUSNQiWSc3vlh2YmUIOgqPywi63PeeQfxsj
/pexuyQGvESLEqveHjg9mrF2ElsYEDIf1JbgbxE3z6MypmlPu5fKAY289TtwazxUQdyUrVPJZbzL
GbZFx2KQ8/LPy50e2A+xKAJshzAmbwYQIJiao1fj598sFmIQ5oeNTNJA4mzmPagmqoOU9hpSS8Az
QFpe7tBoCo4LW849lkvn0G4eBKrGQnz0h94B4Z3jc1HoO1Tcqoy9lcSTxC5SrnGyieBT6q3MQWZU
v7uZQ2+cj6Zl/M6nN9j+U3sL0A2D+5zRPmv+KmyoRP4DBNgxG8JfKuCgcDLuyDcKcVTA0oJVixps
qB/H9ryrgZjixZKMhgVo/2NgkwWjs8ttA0FQV5whlKUKQMcmd5DOqqzC3IgDKJnpo+H/UDkgVa3K
7KadZk6cc7mNN8iKhi93NsbJD7pzEr/jn6f+FcRU/DHC5v0RIg5BjmjyV/3UjRsK86f0ZjOc4zBF
hq+UZqiuR30iJ3psIr3o37sYjJVtQc9oyPUINhUXsQOwo6K+olBvOLKWPGkFV5UFaMYttYaFs5g6
F3cvIgEGjNQ+DY70sqEajT5hMo0l7qKNqxgwSRVpzUJk+rdbADpoM69D11Tvi5nHRZ3BijR4QXnG
az2F4gT0ne+s+5e24PffizmjTKc1762Gp1spo7LPe6zSa5Zfp2Qo1sfCFZQLnFPw8UwJbWiuEIx9
YS6yzvI0yPkhBlJkXM5iMwhzBqW35PGUZug3s6uaZHy4LoeOhP+lV7vWQtjqyuavBpyiHcoe1prT
89DVFH2dflSNsDo3PVhrlFQTZXiAn5x/3nqfUOgLyCueFlAJzNYFwOOrptM1bKErMHLU9YRFDEMp
kNypNeuJPADV+4/kRlRDP7vl2NlrIrdEqWTAQtxqysH6SZ0YRheXszL0EWPYsEwpTroBqHCRlrTV
3hksB/aMaqqzwZmMVGjivx33Od28sz54r+TSoTAn7rCu2FJ6DmfnmZfKYo5eoMRZPEimzN7mzivx
uSTFEYgDMGjZDNYTlR2XRBz+cl4Arav7oDRWDOMMkCRUme+N7MGgK01TL5Pc/DrjH8/1tLWtFi9d
QbWCJxtAq1g4v1Qz4c+zOHyf4BrtlYSo2xgacgjyV1dtXMuW8R3Zea7DpPiE2ptDP18FrVzM86Cg
JoWBOnBO1/dKut7pPvKe3S6bSYRR25xutKjiHdutqPSf3IhtG0CXa9JEHvTyvjGgzd+X2lWvHliW
JRI3Bn6G+0i004KmL83qel+y4Tu8RfydNqbgI+5REpoKb1cxgn8EYMPug3gcb9ekyFLzW9+q1928
K9pXU4e1MCZ6K771J4PCqc66u/VIg2q4v/JJmGZT+0qdK0xV23DhwCHFuLSdR98b6vN14ZJSPLJt
NreC+ALxu5uRAK2eziuxAnK8E9Qty3yFYE5s0rFkiObDBzl+sfEbAgmZUd96GFeJoSnLxsL71s/f
djBr5NXWIstCRWCN2N5D31ZR6gDa4EjBN9VYUUKrXiodxhselwkvbGQDfhIKQZ1vLc0k3MzU70on
u/kpN+BSP91ZFyMvMTFjFCE9YFN1gLrjsm6IqEW0u39zhjKMIYTgjZepTJMac348QpSUP+DytssT
pukTUBPW7wgNKV1ZkGe94HgWL7DEwN27M9rwC5XD290TK4lQEhEl7zY4WpRKdNoTQ6dPQ6lM2Ww1
WcNvkdIBWkiysCE2TixjvY+RFwBNzOkL39fvO+gJn4PHjAuK6VSv72lC7kObLpaivyeenmTIVL12
uICYAPaaTK7t4hmpmbqCjWV1PldNhPFAd4V7GXDMk+DliiIN6W4pcoLf65AP1PGtghlgGCL20g1L
xQL51Q1IdACRXkBmNhM4R1VkrtSyyeqgH2rhDvic/cisYmPjFcrgOfxVcObWtRuaazsr2Cc7eZpX
KbSDL+j3w4QmRMHskNcRVaAb7hpsdpQdgNGR30+UKHTNge/FcP+Dwf2gjQ/rjABI3i84ZSOAbva7
LrDJ5ltmkUW2hbNdkBe+jC/CT3RfL65A8VyZOfDbMUqiBeTofQp91MxAtRrNbZW0B80q9cmq+XjH
D2zrIzEaTiXPtIxvFnEd1CC096AorAZTDACZWUMNXjeLZK3GxgcVX8VbNAR5fzctJB+wXv1FKSvI
NsVUA9snuDV0Q6gtjQTKdYYOWZT7yaaEiYTe8d/zQ+ZcNnJO8LY1uRsyxoPNxremwjoaSTqTvNfH
OTQzirB8GAh4ApyEvVbBDW5YrbaRCxbE5gs0yOpCke4z07Qf/9p4DOG50jBVO+o84dt3CCdz3zl/
Q0DaIzgDw6jDvY2Nuou+E3uBeMgClPPCriSO5sQo7LiSUWu1JkhZuOaWJCYcfDtdnoSGGNoULqJW
YT2zLvo+J7OXDbCENenGJ/hO77/DJr36WarfZ9uwu6scocgU2Ljgj3q/T8oQ2LQYu94PQ4LsLfYO
S4B8GC1C9IQT7TkZlNUVLQa9rb+xzKkGaOWgh0+tGWRJ0+JN8zwXNPG/C7v19DGUp16OcFnpoX3f
4imBsel/i/jWYPbfqShV+KqALm3U7Rnjg8bki5kyoFRE1JzG6kCj7wx0gYQ2U0e+rqmXibaZZrTH
m5KUa9A7SSkRMTKAwVsBKC9FZSg3qHSvHGxbUIVESS2cKSVZBtXhnq15ICa3Rjo4pRuIK0aanu87
/zhQN066xO/EaX5mi1iKBBOoSfND/Dmc5y7Ltan3QcUHSo2qNB2Ssx+R5vcWKJq3+tIGReToePQA
hgRjvOPpCoLBcCScC6Lo91XPs0O5O41A3a/tQB2BUa222vITJSq5pVpBcVlylYgjd+BUlWrBIQJx
Qci6lIb4laKoUdJtuskKeGE07EyMw3pA9C7nzsUP3KBk1VqSwfl4A3lQIBhsUFZPM2t7a80TNu89
GRDj2pK3AHEIe/6aYmilKTAFSVPDeg0P0DZkobMiO1rxLyDpJy4MlPA1ml1mHHvqnJPer7BCXfHM
aFQcYNVsWNZg7LcV7J/0DItF3cJvZHCe3NFVlgIZmMVzWaeHXFBE9AWqAyKAUHDy1qHkFg6XuQMF
2HX5P9bLzAWWC692Me7e2opSnp3Jk4uHlLITt+1gC3z5eNKFKFh1oLtDekhJNBcBsLN7VGtfY74p
EmEeOMgCidMA26PIa7xsLszgRm5CEHd04Ye37qRTUcBK28sQOaVmmsRcsX7jYVzABLoJ/1uAUC5U
FDJAZnCY4vWELiL8ZrEyz/1pGl2qwrhlOdYF9kJUf1uXwGX9MvT0SaqCmP4vD9Px77gUlUVA0Kda
4Gc0XtUwuRzZsj8VZnQ2T2eLNLbeVDe377bZuRtPuLbHM30Uir5AC68XU1vZP3UlY7DUTsb/Y2dH
Y5RI9WmCpCd3s9oHBkqaMmWXS5D0dmdZZsoAvguv+89aE7zcANochrr9iD8TswbWd+22gDFwgr/i
aytde/8S2Cjq1/jAt1jmT+4mT9LsUEGG3DvO7H0N8tU6rgCIPtbYHHES8bYyaKyrI24AMMfaJFqo
N/WwywqYbs1I5rTGA5tp1FoTrL/pYEuqyCvyoM56MlPj0lhy0BZeK+LmN+DaSVRjYiPsF2wsLs/c
HKyytImIOCVLwQ7VTRMaa46258PxApkBSSXHmU80EjbGhQ8rzr+0VL4vTwlqwUMQLu6b3l1KypXf
90N7xXUFznA2VIPRMUS60LSEmg3CKPvzrZBpgrt0n59eQ7XgxwlYVWcvrG9KCn3t4MS61LXBSQwg
ezowZXiiSYeexO+UJCpuH5PzXcBSXXm9hQ1Ga+tm7Dk0cYob0FLNPZrrUheBvNEN6YW1yxAXuTSV
hXh57BPcqefN9uLixyxkuqk8NppOVUczjY+Dm4ev+FcpIokrHIg3K7zewPvh3NuHJJgDRG/dbdMx
ptuhTKONhaP3JwXUlyOxHP/Hr7orRuotdJzusmUqK6sTUOUwwepIJKyOhy34JEO9/SW7as+iYojL
TPVsZIWk/3OoDFqEZ70r8Ve6DcVGXKekAno7vbVMmOgqyggtWcif1T6/LKMxq/0J3Ga+OiOJ+FDx
tC18BrLFIXgkx83n/IPIlrB4S75cXs+z26AF3YzIDRkuwHwGmgKyU2V2ccWvlDpsrcDyUlsSbGWN
zDu5EvOHltvmW2AoyjEBG8UnfbZ7RkgW+nvyHM8iq/fUpaKxmM7rOfIJUB4cdbYZRk2Aq1vSQGok
j7KNfqmtOWrHnTTfdlo++BeGhOwltB5Eczd9K4ipDnztAohO32PSIvj61OzMHnwvUWlP3f9bFAuy
oit2jlr8ypGF9gpSbPz6AkVcgLb7BzfQwErgO/baYKVAzXDUbWqBFAnOQidk1xySl1435Udvohpd
Bt/oOtbG84vBAo3GsZ7O4TWaVmBZyhjcDw9KfpfuVX2HqDK3WxWP8LQwkUSAlHjzzz/EsKhn9czn
IPw75E8lMz1TnFUTTA18hOJHr7AVwy/zsS88YZH4WsMnmHcGzmdxuyu84h96ip+9tWhQPIyUfuH3
L57ljk4zbojW6PS5qmQZqBudp13OGMta2WUR2R9Hv2WwI4h5+hkiA4ilHpa6aDrkqWkUyqVemsRD
bTkA8cQMfGoiYC8exsKu0D0WzKUWqY5UGKG3Nnk/2BNUSdZsxibnKsxs1P7st4ak+QyKad+FHoZ4
JuAggbDcyzW+V3MlvYBx9e8pYEoG1DkTzbkmMFd9C8VBzoI8BryqD4KuuChfd2sZ6ddNyfoiDhb+
Aoo/TFYD+/ztXz8NqNBul4pubDOvecb1BX4DLsBWQd31uoq+fHqyEWywROV3XyW1KTtbFzsJ3Cpg
+rMBGUXF9zq/G/x8OieXdzNe8/DAOxM26zS1poQm0RmnS8wVv/MTSNKQei0Da7CT46WwMfWrGqXZ
U4DLjwAQVQAuwTMf5m55l/aAc/XbxqBmYODpnr//8bPHezNr9kdvzHZG7lcNiOuDFAb2c2Apjo4n
fiL1mAqseTyrE3BKml+HzsFYQEJN7Dl0J9wGe42vgzzjt0f0OHfArbyA+h4ZJ8wpec1YUcsLvYNE
lDa8uCeePetBnsU1gLqbOc2tRxlKzUYvz3x3P0d0tXXlGinEansihP+VfMvrGYzWjSTV8rGjul2F
zu8L1H8xdmIsJ+PWyAsdpemlUtEZ5JCYucUrIz1pvauSyU8EiPXFsaq2hZyx0UbxqmFX2DFdY19P
iMDyxmboE4rj9ovWwiT1rtDnUur75TCFHA5qvVvIJ+J4ErijqpBRKrePYAUXHAyId+GFJMqx0YXe
a61o09YSK55DBuN2xyvL/LvW8u22kQ5Yhl20a93mgUHs0m4tleOgcpWprYitcOLuIByH0p37GXrf
QsUFB/X68+BXyQYL4LScn7Y8zUd56ccLJsL1nleX0X1GuVlgAfdRkPMTany4B07nQgJkzlQQTf73
1M8kHQqghcfJUlics6t4WDYJYoiQISaXxnz9S9vLVeHezkIrZggw+ynwnnpbJtpofEwvOfcpYnTL
UXz85COUOFwk7+KLdeXg6F30KK8HMYmrBYJdj6gfhfhAyHb2NIhYb33e3kkNOuKTeDVRmViBz/LS
eDyZq66NuUPpMWS6Mtp4M84R8tyJnMGWS7c4MKlVwbCRlCvlHgvYx2yWS4btmiGhW3uxEjtTqwgI
OuShDf8pbAWfOMvA3EuZjfB86FRDgeNp9fTAyMSLHkQ9OLaDHcyu3uR++h/oANoBuJjGnLy6hEL3
k2ADOAKIHsfAIgljoAaGOjqQEVi4qPLvBXJc4ngjaAQDmj/xGR8vtV0mgQc/2J4FXDmqB22Dn4ga
ZIVxfZRYdZzHAPvsebrhBM3d+a3VNUQaJGihppjG29ExPY6mlU5Pv5smZShP8I+jz5YRXbHFjZjD
yywRKPHVuzfJNAiAnBSJ9oJB6pY1635MF5qH/VKoKZ6N2C5X+teY/ucnJq2SXKCqyuQpix2hFsLj
N7P6GdKxoj96n//R6Mf9v0YDSWnOiTBr+iqXmcLNmcadDHR62dkVCXFYrbDHateiBTWwWC0CVcQ3
w7pWtnpmjGX2TtyGSSmZ8TF2EAML9XJVwLfF9SxIVcOi5ddUFc3Gc7yauIjCqB2uH+48XQ+AEqBd
wdSgqpnM67/jNHP5yemfpuuMwHv/IM+TqdG1oT3f79dMpxC8pdooEeD9kiaCsHwi+ionq/w3z+Gd
6WIOCCLOZW5Ws+DKdw6keGyxPSt8x+VE+orIWcy1RHxejWm3FyGa7rOELZ9GXvcKXiEG4taz0taK
atb+XTbprtDU/Vob7DVX/U0a3A5iIsQZrN2zNJoslzK+VDOTNLqNS0I84sa6fo3jUMULX/yISmIh
4+19JuON9bF1VRRrYiwveMdOaysxHcL5IRRrG3tnqw7DZR8oQzdDH0n0tGk61lkGNbunQfWrdYUe
fc2S+s79+atyp+WXHmwE2zMhBnhMxIhpmX0P3hMgGcXEFCIiyfZ5SDHR1za9E+CT6bBu+7U+ITOu
WDKpD7BBLDoW/J9UFXEXJtnNUxlf80SoDFugbeqsogCyz8TId2AYo7W7JtXymthhMAvnPfEwAOGU
2fw7UzgA6V65q1wcVhyXHGpWUbPZWhbKhBRpZXKRuugn2zB4HuaUe+0lViA4w4yREeFDVnobWHDs
Igy1c9dzTTcrjt3U6WPeE8BSMWH7jQx9I69OL+IlnDHcEa8E+sgXMNgggeP78Do6T6LDrq2NeYZb
ckMTA5nEEdtvVdlBKcebZIDW3oIJ4X26zuZ5OOxIRxaSPtQrWTvxgSxKaXsedp1tDoS5wHNSKccv
dvTW53Z/PHGzPJfCkMGfwN68DPP8DVXAHh3xWbmiH3Fnr9HSMccs8GfoiYJ10f6OTmuQbyCIX54R
jBtpinzzuHJ+C8CZ+sbGuwL+51MO+DtyP+4YSEft6uHL43mMYDaXc4Nj34r0ve4XaEtlhX83i9Vn
NLERYnrV1iMZUohuWNUCzV4fecd+7a3G6DkZOnlVISzmMARNNVNAb26gt99U/07X1pnx60B5UUw0
It8w9aTrkw8f7MYt041pZio+dXl5epAfioWPU5oQilunmiXIgAKKbTKHCTGCCrLuxzZS4X2xxL2H
z5vEDsqSpQhsROwOvXSZNoFiGIQFCywbyyXmgNnU0roAr5GckGrvziG7VimsQkduhrVTtc92+Hse
SKH/UV+ZJ6r0lMonFtftl9yoA1uDGNySrASUR3hdLziSvyLpoFjJ7Hz0jeDPfUeaH58n0bbsQ/tX
dZSYY+HcC563pprAeA2B3aao2P+e9q+5ru7Fw3ZTt/MQAoW5hy+u40DsluM9DtQMBz0911pjM9wQ
/tKBpEol32VRTdMqORzioku+49oxiK58BKs39u2/HEo88r8GRVjRt4I2mSaYXc1aVXybBoWnHQxt
lx2rFK/H8p/LVESEarRZ1SfRdWVLfn61FyP3nPRzKCbnuqKvFnnKtsrTt6CMsI1fpmSkQqczH+6s
9g1b4D/R1vW/yhZXr1EvYUNfdIzbK5pY4y30BqNT0DOfbZ/mJFLB1L2GVVul7afd9EPNuQhR97zY
tLyVTw4gBfMndofnHNLoS3WcIZDLhI5BH4S2ga1tnQFkGzCCuGdcgjsTB42OyoLP8PkcJVghBgTC
EHPvlHU2Rriw1RIYEAYclsNq1a+Ce7HQNEj0t5GGGO3Zj26bM2y42aRrxDMS1dCSUPU/P1ecgFxj
ANChbIcGQdVgQbQs3deGplp8abqyNNv0OwzB/xHSSnnIlqvK7u0FFp3CZGgUMXaML95Je/1Tp1na
aMeGThvZzkemR0nLqIq3cV5O68fqD7Bx1sUbHXtl892+sR5vC2Tvy4jmNQ2t1D9yi7RDIuInu8Jf
d4K89KkzuWURC4jqccvTP9i3nKYmPklxV4oaG7OXxBauHN+qBdShWC+DslyJNElGCsP3fjznWz4m
lvBleVZU3qJi8x6+XuM5+uWNCum4Pxt/FUCfwDF6s3QauYj7biNCos2Pnias655ihzBii7xhyi9a
elW49U5dHo2DGqKOI6rlOdCVWG4svdVtmyxY3DZv8CKdNww+B3fMTBW2lPpaUwgTgIA+TTLjfePM
x/Xyk+5zLSjyub603K0imTQ0ySYhG9OZknTthtWK5mYJZZq7VyHzx5adptXHdQTfYaaB8SI0Mq2t
vP1j80QWMaohUf9JYjHNp9bNeImfOasvNoxKw4kbBHHkraRqARqJL+uiktIDE8Mx1ZYRlFKMuY4j
L2LTx/8ITt5J1+Wol746p/Qn1JBadDmSDAe37xYVxCdzKY6cYUyeAuEOCeJVlbY9iM1Q1b68xfGW
H1awgqquAY61rN+AwEbP9oYLBVavVVqXuhok/IutHrYz4uWVT9qIJlcph8Vzb5FWSD8YeOzVXQVf
IFx1Lz4J30v9wVs2wteuag76XebgdQTincm/Z+ZWuWKSYqvIMGzn4TiiE8PYsnB8U8bAWiLH300y
mqnVusRsumuVmA+qkKLTmJpx0SjFwigL+wxMAFIYshuC3oaNgV3xxXWqslm8lIXt4Ypv7EGR+JBo
m88Ijb04kwT74lIViswYNh79V0pJvgpQfXF77SQysPifpIU46cg4dOSGnC9GV0DjjVEwwvbH5WGo
xuh1lEmrE5iuMmQ1BSKvvx2BwNLW/ioiVyhExFOnph2E113Fhj2XajAprv/UOSqvctYxFeOBintl
xhQZ4RDoKXLoQnukKDim9vK224B8NMVAOO5m34BRfYZjGTZhieaaICTQ4xw/ps086tnIE+jZZ7tT
vqcSsPgHodjEQRDL7YxObu79NAWBNr2rCB1z4pgasokrn5I8ti9Txc39D16mhShv+0MI2bhl1b3R
4WveWQTsQ/cL5fPqwrFHVQG5CU01RdB/qcjws0ck9aSheSVkfhbnVh4LfXEv0yYgpyPgkmvE4cWo
J9BjgI7AdNYH045vHYcdSQoAnLgVkCCDl2Z+tlkJH+UjgvTSj3DEOsjAP0o7zs8e6Qc996e9bdQp
mkYlKUgql7LMpNac+9+29xLuXPzUINNoNYZNfOIL5Dp18TXZC4IK8KUn08ktAnVMTgiUws7DlrrY
5/mPo6kGK49APuSsy1Do7Oy0QEsg5yO7famR4gXx49NzH10aL14UXrcKqESmGdan34owYLNOgecV
T58JpKh/OYnbaXKakNsviouyzI3wIho01AUkQaoVddUXTPVKvTHSPj6LXz5DyIv4fDI7DlqDMJtu
jpBbzWRE81DrSYAUMBwd5lrEAGPcWFnX5tehret3hudPoxBhXZSUOod5F0BWuUDK6RkW36thh2JJ
5R8GHm2bekQtjqUGJJvJ79NwCBqHrJHaL9Om0kr2NoZikCyVdxVPRPDk5xac7SnyHJAkV/ACCo7W
fA8lbbGWHv/UBTxVet5BTv3FUaqqDvZCuuImXo9ERyD/SFVtrIfU4wAe9YPM7nLNi2Q+88DIN0Kp
kY9yif1fd7Mz75PmxKQfrGFXq5AdMv/yVO8KiYTomWDEaHpE0omhtLccYS7KFvYxYozPnpmsF9IT
zSNytLxAse1EYafKPdNzxnN8KkIvB7F63HKvrslAxGZOFRCr2ncb6HrtqUY7YnYpSobaiLzThRbs
hrK39UJunxgCl8xwiY/cBeOcfwLvkkDZaC3qr4+Y18wGsvCDyl6wGcEV/VyfCjQwW2eUgvXmasgN
wLnGvKfc6CFxqPmSUTxTeuMlTua8htlg/1bfGT8PbG+p86lrSqujz13XA+h4SCBe7opR+2Em4PYh
nAaBZBTVrKdkX2oaPo7c0dToZYcR1U4F7kkTUdMaXlUgRm5sra1AirciCq70IL5Drq/B0z0iP51K
XzNjrxwmnsn6KTLtbNNOXSN7h4/vAqdzGXCVXqQGNKxUTssYUz/D8Yf8MRKYhpDtcyDw2fooAwhG
+eVc0vpPQA3WoCJPSFD6cQkPtEj1ipT0L+fkmYogKhbEzuvbT1PIhG888CT44u2mjFgCsigOZOYG
KmGlI/hseEjoRhNwRbYGglvtcyepRqGwU2qWv/JKR7nC2SFkb9nztmJ4+ahvfHaZ9WPWntZFGcYr
RpLboS/7mZ36Vo7b20l4/DuhUdHo46n0+PX2zufB7M7SbWndIeBIneihIMW4Gqx8skvquXr11R0J
4iIk33PtqaiC9vU37BFfpXibqbCk3G9V8FjC/fgeHKhwGjtgpI+Z+Tz/gD4e6lK+S095n4dQYmdJ
pWpDrecG/zd4lK2OMLQUiADW7SleCYQRqcttL6OiA6lJXF9g4SeW8qRsAEa7FPh7ARJFB61E6L+Z
oNXa54SEKXqpibj65GA7fBLA+uDw+XdDSlFkC7/4ysKp6Mc7WR3oX+fkM8WHfi0FnrsU7plzEVVY
GaWEv6wbsf9MMMnpQPZnuHYm/f5qm3jeaIIRax6T4MgAskacZZORE8i9EHfBkIwU3fOarpUiF/TA
MmO4bipJ0uiVMeF4wUhDw5RDuOjkbM/tvf2sW5kFn3I0jua4Mtwd5kpKWPtOUlH8aooC9LhLCh7v
pJKLcdJUwGIX72T3p0c1vc2bTT5853yi/3ncLPuoQwRwt6rMkoAZhKI3sIsnWqe2utEnZCdTvko6
V4EqSHg0uf0Z0Lh+pSreJzA/fF1p8WCzWJ89T8QzSrUWh7IynWtDhUmTipIvMR7Vj5bNtXVHX/GS
qRrckG68MPc+y5ZGBf+Yi0DUHpiYZO5Krcc7zoHx8EI2450nF84esewcd24pVuvxKrwI1jNKKrP6
wlqWbCOY10YI2qDNECEUv29fjdriTdQ97mINzdggd/WzadQ6yRHScKD5N/HUcsX+paBh0l4t1xK7
b67AvYXZoA+7OZsBGP7LKhIxHb9QPOiSdZDxXQeFFPUkWxZUIFmzMdbUpb7cNkm7qz4xPp0QWMqG
D72ipjP4dXe4VPmUd9uvUFsxR1Nrjg4K3eOU6NTvmndQ5x3qaEZ7gxRU5LU50Vqqdh+hUB+GsbTY
s/2u9avVyZONoqPO9jpB+29Cj7MwCnERt9OmVM7pT5ScSaXZq8Zs0JeaE7zCLn093GGKL9V0dc0s
ia4WKEaJYZgDSzLEGK8btOlXtZQy9iL0g6swCrQr6uj8oqELT2WWwWQMbjEJDy2ReUngf9H1D0dY
Bvzw9wnpTfx2eBqrjkgFG86eLfUS1Xe4MWdnKqWdDi5JnO8e+MmS4Ov9nE8jM7ibO+MkuaF07Hwe
rVy7zmbY2dEdi2qR8+6hLLrMyv5GSol5j0/PDh7R64HZ6se20Nj4MYiD6f0qOG3KO3xECa3QY3MT
BldjaLQxS//gDhSjlqM+EPm4rhgC6tiF7uJf8JVQQNYkyfDQuAv8ad1G8luzgVGyJp4ML7eCnvBa
wsbdmQ6zIYbsQA4Oa4yTT7ObXNSjMNvNwjep7q+i1oLjbewLX7xBS7TgNzHc9MF7EPcEifV40FOV
SYlFLC9hlhq4LFSjfN/C8t6hYahRBthb8+yr8G2tCyczdO8kK7t82Ljwul0bQG8sDRxQktlvph/h
waGsJ2rxqz0Zn4IVhDI8N0kAsVYN7PqDqr0pYidhmBlAkZojOD2gcXBVyoKyH2RA9SzlVA+hj4m/
9RN6+c2Zh7E7xGflCAv6fbpITdRChoezy+xw4D+5c9pAxMTgRvtpCGsOwYjgyqOCrdMwNIk4Rruj
KGlZbhp3jSuOpFmEwRUWyaH1D9aLXTKQ8yio60UfgZgawu6cnX/XEOUlloas6e+WL9T5cYQfb74U
ifBfNkKCoY81XMmRacUGzSY67serDFYQxLKJjdGwXnuEABXZcHnUQl9QSfk7Fb+tujMj7P3a/Y9+
VBzCdisezrWCgx/W3yX6LmL4j9bvlnmLAjjZAwcNdHa9q8VW0T5OxzUtn/WJ/YdcQImT07cESCOb
hqgpFWlbKwvYGGGPXGeI7sAwhgdVBviTf0zh0K+WtGDa8QOsomvgezyv53ieO/tN+/kJPL1LY3Fc
+HaHYfFT2dNQlUFlF7fynqrdZl0b7XLqjyG4cwwbyyTRl/mZL+d/2I9pnuojhUNIFQconHIMHPct
/6OwaQizOIjFFLbEhgHs7+TY3c1qn9WBqOKX6hCupOjpbaHzlWBpwy1K3MeLy2uG5vgGZbhwTndx
X72P10ZwiBohCQ5tj73A4rZB+EVsRYUPRHmJurkH7wh/2zRw9WTHhQcaaVJz5jnUU8py97At/gO4
8Waj9uv04/QYsHRGQHsz2BNfI4ieApczaJOK4SewxIH/IuIe0FGwoEWIDEG0iGZpPk6uuuuZ6Jpw
eefpeNt4FhK1sNELseORzEqT4qEnW2epJ5p6M/YxFbhqYpXUrx4Q3Gb94e1Ypt2ty3684Cni0oCG
mOQwwfr8br+dQGnLhPkZOjaLIwjc/b9Mj4bfF83Y28snv3OI5jsQEVdzru4uFbZmL0yoKC0RDlye
d8aqguhX3IDVN6vNJwnqmsxkbcNS3QcCEyYMjpFHatkz+6leyE7MYd2W/cUHsL3jqTfqt9UBQA6T
RIUdtqY9hKl69ALRLAMFBJ3oM0lFt3NPK3D6qL4srFGX/3pjycH2vCVqikEx61KNWPv3o9bWzFDo
Mw4e9B0CnqKUB5bKJgm+5EgTF5/nlh9AaBK33PeU+ZZD38UP9sqLu8HMN/9QIukv+lXYKurpOdWQ
6fAOoNxu4XQ8Oc6GdEEV7TLX83Y+EVwE/lCqTTVtTYLMXbIJgpGCFFYxMLpogvc4tLgprJBkzB+u
p5Hve1Y4xLQypsYCPPtp+hDfUPe8KuZ8sEVdCk6TMBYPT0cNnxeDMQA+LO5alc9oy1E6ypsUOCR8
Tpunst2ntsBK+9AY50NDb4OvVYt9javZmNuXlYV6RSR/grHSHzJfG2o8sNN6023dPiO4qOkmTnAD
L+PHZPmfzK2ETXLwm5sRUU60qmZ9Vk2lIYOSqoL3gxw1OpB5iAiTiPHU34gxFiYUBRAp7cBwjqod
LovseZUxndVwPp5fq6j5UtNiXvo05gxHJ7cNybxlwOC+Svcr7lgCy2N4Y9RtyX5vrDrTT5POWjyG
9mJfafDvw+tdjB/5OQs43JBtx8tcM6GN+7Qr4uWuOhvpdcvsFbPUQs1zvxIhikph0qnUwXv09JN3
xdVM9TYSHHk5YFAVvHvl3qqGaaZySSZJ8LeGl28DdTrGlJJxBVec+TmcdrNSlluPjzg067gNqr9X
ni0TYQBfD5J42P17yVqe6VrPtL47qUGgOl7WtUIKgunDorJP8eROBGB4Sila+dhPHm+p/S8+5wyy
Xfk4rH7+VRReUq/1vbOXfCJ+NAj8aU7Hjyhounlg2MC/8QCmNijef0pfqnSXsrhiSnmZrHhapHfn
CGryEVfs7LsWNbjz13l2B8X9DboXf5n+SV/BVjabPAe8ysxG2ITfdDnnHZ08UcUMmGvgCMDOxxBH
xLjdoty2dS3WGfdfqCebD5361wHjhGaMgYuGtxJDE3iNL8nn6cOKXE5mVXQzGq2xJ/i/LtbM9Z5u
BeGpiIV6b9ZZ0Biv2QpBHmPZ/MuVTuLKXi82z4eIE4oPZeuXGMnCPv4AdZUDeSAgOIxgfY2c/krk
6luETq9L9H7oOzL7uwJW12F8reQgHqe3uK4EHOtqVsPn0UOGWjSbKRN0c/FdAS0yB0c9KcEXdjLf
gV4s410T7EISuRSGsp6h/E8Or9Py+6Yxs3sTIoYarIKbQfBzhaK6Vm/2/riKBvXPq+hMsc7PYxDa
+tBJ+TAZuWlhhY7lq/zhv57uCE3vY041o5ZE4iuBE+IuoHvK4eDgvPymhtVlh0/nKfm5pxi2gFAm
fC1tZoB2W3qO8XHZw8XS/8Yq4TKBeARo5dFVJaFiCauUDAAvw3X3Wk35hl3NOpGvB7fd2jY+etmN
y5f3ScRerhwXlpNaJYc0Z+R/JUTfNs4akD6xN5dbx6m2SM1juhUqxmWZQTjuoU3mComECLYytJCI
B6Qw18kqLYC6T9tcGihbIXdrZXf0eDhf7kyJfDHMb8faSDmCR/TVgOaQX4bujK8e2u4bseG1Z/oq
NiNGL4sVzC7viqQSDlqdmbUc5JkdaaW9SuUMyKssUWO0wMI6wVDipK/Lx7bG8DEtRKzISEjHP8ja
pIRKjPB58hwQ08NlNu3937jIMuZpfU0crUNZ/6sjLoLmpPfWNiqYBCrSbCZH9CZ576o9MS0FH0vl
7V/D9gMxPCTKfNXT8Bt6rP/DQd0VrZYoP065RKYfkFp9R/bQ/wFSQJI8jJVFGwWyH25c3tw+4tvL
T6A3JTPd4F8qErhdVh21420zeKUTd9YGkdhy2+xUZ6qLqFPARDDboViopf8pcSzmp1DPi89UbB8t
VrYF0hQQSC3hmAHqR7YZKdlyphSxi8NYgTNWNQHW1KwuVSUQnKzGPf++BMDvt/1xCWDitC8qGTt3
aQfSInCrW5VNjyr5zLa6vJCXoGJi+uzCFc+gbDA592cd4VZoQ0E17VBsiHd6f4bbtCsPqsmMmWJ+
pj+5KdzrAypRouTA7uep8vKTNYT4navPfaMEUamZKNppXWMtcFe4H0fArpzU182L/vms82ALiLjA
EcLhHfzmz7kjMYX5nH0cSp7v9lhIyqVPF/dOPdlyylQL7FC4LYVyQspqQdlFmUiIL7J6C0jWXB/i
jQfHdsjAjOQVHQEzjclqLsBv5U/QLTqz8OvRLmLQmqtvcaLV9E1fqTi0cbptJfwBLSTHy7b2Cl+K
y8/wpjLIgnVvtcrslEmAvIadIBqMonh+16xBuoYl1CBnEFSCxIhcGGZ6c26Zsz+MjwC+T0jRvQSZ
SKxhsompG6TieroRTXuxi0Xhv4x/V+ky7e6YDZxZM+OUCtMuYoyXNuhWNDOFfTWapu4m+kKYjq5D
b16ChMJuIie/NgP4WMKOdDYWo5epNeFoy9yxPgj/b1w/6d6XZIL0xF6eIj6b4vPtG9A9lsIlr/Ly
y3j0gSY9SsCPm7SBkxPkbyr63A3TzAsBHVCxH4H+d0PkFI40hfEgZfCgAw7CWclaTkt5zKptGKz4
m204Fl6yTqELTw4LPeFFamFrQDi31gGKNzll1udLcKEi21HLB4J2YQSIMhPTIz5F5zLWOh9PI7j7
5v8k6xB51FpwfR1GW/X7O0bpTBk2JFsWAhcWXfzlqCfcU1cHiBYbdXlpJ6W0/I8siBNxC7/d8ubL
9pYHrpUkxj05w43ukfxw+vea2bG8ssb/pvTgPinnpUbrhTFBfW6DbwpjfK5+OSLIBU1JZM9c0Ttw
SYFwxRe01eFmllGlfRWg2W2NrscdJBGsvgp+fqfg7OKZGdbW5jYX9NdL99pPt0prPThyrF8yX4YM
Cj155giFoWgtJF81/PMySq5Vji48vY6Lks8rh8XjQADAa4N9RpeUWNdIY/eDOtNz7KRVAEj01a2t
5Po4D9wxICEdtxs3LKOakaDUbZh5BbTFHXPhJSqmqfPlxLyhQ064y8KKmWHfPfAaiwYPMwckTxML
BuvQNUO6EMPuhZhm3kjP4hAHtUjz/L2sB8JSSq2SOyr5R/2dTZaJA8agXVfMJk7MxhztGezm6d6i
o2l+/HmGKxtRABQIkQSPyNlJz7cTCeh5AqbFSpwSASEXZUnP8ogEJTNJ3pphZ5zAWCoYFWkTmwBo
C2dBSXMeotb5R1C6IqPFK2t074USFKBhvAR2XvE9r8LwCejMsJMmKCsd1kYsYqyvf0SDzc3+7ue9
XphFdcDtyLbuirTVlKa6uUA5Z3FOMyfvOJH8M+jMzMiKDr91akNJp86sq6C3r8jVp3rlO+iHAykz
NjE6wj5eThCCn0xkB03/yxA/LwEUkDsBwbHqoRl6OCUXHVLt53WVIeUaUYIBpwjaxDKO48P0/L5G
kiaBbMz5jyW1nOF+zKEIOzQu2jEDwoUHerPQq3o15XaDbsHpHGHWrsfZoWK9YC4lKFSnYWNqTWyG
Gg4ZE5CkN0SUraN42T6MpJrjifD/gXXM4EQE/+Y6dIchiItzkh3MeYcohxP2hWRJGLAQsgfBg13z
Y8Oo0ROpRd+P5wOzCNZzC1Byk62t3bGBHaT846docI1Vbb8tdSZeYlb4Am6DKGN4WCeHdNaj9o4L
nymmRG0aek5tkdyyjULqOmb7rBBsA40UNareP7IAiavOz+Ae3pwwr3NT9PzKUkggjdT1zD/yay+n
hxUfim7CZZUgUNoo9Wal0C/wp//5XwcJeN7u0dtRII6dk75jQzn1SLrobQL+NDW82dlRH4WIWDdT
STf36P+4266q6OUdTeZOwtZuDiJnW8pofYtfpXxMPdv7t1coqNgo3DfkFLbpMuTotNyLJauHBKPD
Ptnwpt1PoWWx4VdDLJmVBqJL/QLcti1GNJMNI3ALRymLT2ceMIaLcrZfxpm0LLSZUbfRjtfMGKmA
vF0PBJZT3MPvZCKZt49uYZ0diHD6PvYJFusz/sIvRsnqe/XOaTF0Af1vgHUe298r1xLnMkeol3Po
U7nk5679iTB2tLo+K8PyygbDIgdsA87FaUsYJ/wpYXWUBhKb9aXE3eOJAfUP14LuKbAafzuLdvPD
K3pXT5hCEI2pYzBDT8GMwREkplSTKWLeFvEvnIQeDydnZi6Slr016dj9DTT2kGPRAUa60WO4K6r0
U/tH8TmPmEKNUrqeNHe9K8teDQSkUW5XYLpEQ1zbRHJmxS+xw4P7jphwDs5Dy99orx4yByNBCp2F
xaG8toFWcKr3uervNh6vvZSb7gkUEyQtwZUIahBZqKIxiaRSx02ZCDUe1E6z38Pecg3QDSIQWfvk
b+iWw+q3x2+HU6GFc3P/3uUqOtb7jYBAdSgd3g1uthByuV+pRxtAOkC6nr/p28iDQv5OKLTwwRcP
54s0FImoZQ02gkoEXBIMPWXzlbELNei0BVoKXYQV2F+SRtfXmoEgA/c7smu8sB8l14I7ewwsG/Oa
wnLf0uROsMQ5cETxw8j8hqt/5JgZiZpPkW73XZ9kqahwrY5szbmyvHAEOHHdhB4vcBj0y7bJQ+E9
joM7xg2CgbN44pasTcKnJsICu+0rWa60tQewpmESDZjCpyw6LMvi0FVPlQKq/VphPwuFpW2bolhG
rzclplDum306yClIamJO4lzyQ9ISive+6zQjo6Fa1zxh5usPcoD4SOEyfK2dRR/AweD6OFD4jZfr
pEUF8Pmkd2ZG9VKGWZS8X5Gv1WXv431RxRnEgmSPAWmJU7yZ6sLGYdl2M4jkpXPHIckyQc+KfeMi
7mbdzATyoEU6qOftAmgzAnhX9C/jMcZW4we198OAgEApS5hvegJsmZY0zXtuINnWBYIYfoae2qnW
DE/t/DhJuqb9a1CvXAJquaEF6M5MfApj4YMmzPE/vwnp9/lj/BU3yHrsitHavx9OA/oi+dVhJJe7
/6Y/B25PyfU136uFrfByd+fc3RRqWAFqppjDs51hDDCqlOnNN/3TCJw/eLniIcRzHYhmEtzGn3fR
VcTX/c6HjzOjOHue3Xv0UFfkeLdNuGkk8oEBjtoXxi8Yk2wUKPp3HilnhUL4It1TKidgzRNgoYln
iVZCmEOZ0GpWkgjImUkwUUUpuPvCX/AI3r08RKSXLG6qNJIkcDhY3thURrKw9nt5ggQ0YXwlXtiG
iw9Xe2i/A8d/HMhcOZUoAdOl6M/ZaBBsenkoWBin0EyFYPX2xfY50cnZVgy0Qdue9nD53CDlw8sy
Zge8cUsSWaxw8aWeDy8NoaxGIJnzm7ZqrYokIfEewSacvKGgOLOJQseAQLTFkbHqB8dJGHZ/AXrn
VmCSBmMDyS2mwehVnsmXUiWHOLPjJn2DhbEEwimhpfOup5OPt6yRn2bjRQ1p+L/+PpSbIbKQX1Nn
GzTTOkxuCVCC3wjeH8dky66DsghgrswUdet7RROLpByaKF2I/PXI8F75MQR42AUP0s8ggmp3CC/t
7kqb7O/ncgecjdzeFZM4Mc96ISVsX9DLFaVMCdooLMd58vEef0mQ/ft9AINLNQju0GnokDiwMmt5
UIwHl0IfAKsYLAzCfaUSIjxeTjwh+J9NEhk6UxE18P3OrA7oJI1BpKu3MpOjqyl/uLlSXxMEP0X4
5oOBD54GbUxyDLaMlSGoxh+JPYcWhREgqvJa38lD+ou5VzOe29N34hk4QPJHyJQSKrKrfGJznjKY
T272W+jTeeyLa9IYeoT5nYA04z94AtU6noyz/liZc771KYND3kMgWvPUygTiSvL813yaG/ai9NwR
Q/fbMfrhb7OfyWYg4WqKgeNuHRSH7X3miE5JP/HLRrimR94Tv7mARuXQVu+diNdA2B15CXbmlnPC
kiHZwBlZ1s1vUCz/qvI0QTiCNU7N3oAEkttqEkFuUU1jfATsvuR9f5beHneWXehFQY2VPSqJXTgG
wU/70wQPqsAiFZvF8IXtqCiQiUDTE/CFb7YLXKw7y+6lWYTSq1tJWouP2pbkYHum70TFP160cLwb
VZUTf4fa8RHSN/mFZ2uii/bYiuJ+vV2DQNdWgYYWVb7FGGmmxIL42SAOXUtfJ3EmMcrDufK1WNyR
IYuaX8WKRDzJBbr7m6/KYe19u9F4/h85zD8eHw1rgJV7jLEeYnjTaWrRp2LvVEER7KgurawO/L4m
OP/tG7CGCbfQ4IutQ+mW40Kq6g648h3LRnHBVj8WneA29Pf+l8+YYqwvI2prL5hJMtLmGNxPYLwE
k4FQ1SOXtREgmuvzOotUEOuk+5FseS9VC/6S09ZJ1jrqvxdjVe+SrzHQ+nqxBW7HFHe1aGD+szdN
NQTgwV02/tOMkag+aWVH6FXsn3v1ZdS+cuL4rjQHspQ3q5RLziFVUTL28W0zLEVwm2SbTKRFQ98p
uNcanQwnjLOGdzhVSxiWmSuRULJEmSlMAfbOqvKRrt81K2dULorRpyhMxJZLPTdw1jfxT02xUltl
UaqmbLwH92yBfdqr9oYQI3zCW4svV/A5BYhFdcPZPvT309oV7WsDpnrbnK1ektOVOnSVoGnjGdrc
qAtg106rQiBGFmrIpe4LGYuMJgaSaveS51IqWq/Q7NU4MPploF7Wert+GBB5WrTwZ9ygm6kFTi+z
aXgPdZMH/VQZa6na6xl6JZIr/p8UdUUVK9YLEQqZzYKkwZtRLwZLcqvwgt3tQnMHE7eHlwMEMDep
+sCd+jJet70rcmzWcWIB7GzYFGgGd5QqHvkDEUu2Q3wlVfHPUJ/+mz51kStSeDm0BWmAWRg23wo7
KOaaWdmm+EvD5RQYnXqKNb9lukl3j1p86Qbl8V7LkFCiBEEUfk56SBxrpnct8qnjhEIRhGEFhD+8
olotuoDpU4rk+AwCqIBSUTw4I3r1KJmGYGOPPl3caOKCAiK5LRcEzxAJ/b+ktzm7xJ1oSwfks8Lp
f8kSHzgIR8cOXKhfrOHiB5sW+HtlVYNw8G+DVgqtiu7ZE9EkDV/i3PSeVdKqHAWdcqvanpXL7dph
dcO/oFiA34BPUnQJge2kKZ1xDeK9QSuSF33u206YAWhO4DQxKK0jnj6BNjj+eOpm0RWj0KLq6KkY
wH+g2wymgrGnXEtgkCkiIwLkLiIifQafIyJJ2LLseGMIJ0lGMw6k9YpijfurVQqlVKxeoU6615Z1
biBmADYQVO9XmuOA/eA1B29ChAtkrwaSwbmLXYSAdUB9+/tBU/un41IPQaMGae5PUUNgAR4ZxQ7o
EB15AwR+P5s1pnTO9WSuvnoRzCCMY253Cc4Y9w8Ys38pF7MwX1mUbbjGyEEyrZwPHcmprUd418KO
53lGhH1hyX6fLIfIhZ9/MTMkb7xlSFGR1DwFTek8iYwsL9jlvRvoCTCecry3OOAK6RghdU294Z/o
sUQoLGKE595f/NqnZQuLMnI6cChqg6U/i8Kw5jAkx34NEsRythFQ6+8xFfrLauHBeScb39p0xdCf
acf+VTnvFDNDsKHtS2sGcJH4/1FbmAV/1bblbopZQOBY1k3Nf5d3d2bJofLnvxz3w+9VsdD+AQnx
ikWT0izHqQ0GurLsFfXfl2PLtN3b/NzPXuk8SQ2G8Kd9QavX1ksh931+yEK375cyQN6ZEfQJhZx0
a/jZd0Lx/1j3HkB6bILn1Ob94HFK4LN4XwydUa8xlSzck8aKmEDapPkIDCe5wkaWPwD025CTp5VU
tJfUWFuWXy2t/oh2iwvkxAkxhusyPBgKk0+TqlQ9goCA1ICB6v150UWN8GuLzAcgTa6qLM5yyc2J
MUK9pjCmSCO8KU45Suge89PCw9NdpHsEIJUFN6iOix+U4Zss9ylNpqFSH1czMTXIB+xBa2Wvoyxv
z8L3OUTjIP0ltV++h1hiuqBDuMk3Pwjlyhn0zCb48ZnuOYr82kre0YMUKsS2EdjB7m6NKlBL0MU9
RzkcGKQM/klEQngvEkTmjWw7F3HnnivU5zjJYJUFfSG2S3m+zPLsDyR56cnQgzGy8lsHV38joeKA
77+VV/lL7lS5KTomjiCAi4LM/SrVvR849g0qziqwl2c4g4FBnlAf+5AATpRjc04RgSBbN/3YY2aY
GMcmmu6EUxWxtR7QJPhqpggjD5Y/bYFO1uWvGk6veo/8YyoHfhLgb0w/Gp+3UxiALePe5/N5VoVE
ul2brEWZFy5F7EgcjlyXtNXByYoWr/fO0RphoYmFe1DQYL4zf0m+wyDyQo3RQEYsIUE++eiAdj4V
n2NbMShdNQsNztUbLerjRZ2GbUFPb8aw3KVEWLkg+Vw+V0zynM1WdAOLtt92zuILASNhBCcxPljv
OP4G/ZukpPTW+7Q5xDxN+wk8kMxEaEJpV6qNTE+P9lfqdrpj0qGrI6p1dycKFNhkwCR353ULQCos
9sNAOj5JWRld8LGmvCavCYjQeiFDWQhNVjfCW5WqSYSD4FOiEfG6nWg/eDl9XFdiL72w1xOjymzc
+Q/AzNAKq06y9+zFpV3+apm2xctQPwEr/ZH8Dd1m2s9QiHFc8+Xasg0IblsUmWJSZoOoeqeLYlGv
EliNDv9WPa8GsmRadMLXfpDI4HrBhP03WH6GApO8/sg0i2nxgQlBvntjtxHbuin0Jn8HDlm/7ca9
SS7iMZYSqSxuvsHWYAI0f+gAhPXS0f5Gj88+J3IDzoWm8KV/zY2F7Z1D9xI5s8UK/hH3X0Ct0zMN
pPw7xsw0RiHYn1jpKiq1DZ7pjnP7W3LT3neuB7g2e5IMEa9kS9w21IbUIBEJeiIgl29QW7B9GAk0
mOqCrrKhH4Rssu04tnxapp2vLaLXLyb8ik2hSfQOoQTzZfZvsJ8QMR3hPUgeXYXOf9Hmm6ppoH9Z
L8da4ysBgGAL1k2ATBFgFNP2YjpON1PsbJ+G5PmK2poTjmI+d9Yh36DSXGMc++oDCareUNgh6HHl
zpczAk7tCKqnzW1SlrSrWNuyXSHHXJd6LpDe/0/KLfomD3UQBHIycaWEcBMPxN0sWkeUtAnZF+p9
hthk47Mx38iS+aJK309fxXoQid6H03WpI+PCzAkHAzRnPVEQdUmqN/Md+x+wP3Ke7cdppEIU4EDP
fnHICwQnGiEzftyWKyIOFqFqw0He8QJWFwJ9+6/6FJOohBkvLJ6vZTgZwGCXZuqNKT60BtLD2uth
CqBZhWeSdc82thlK4PdA77cf+P6AoVuUu4gQQ0l0jJiLv5JC48Om7u/j2INnBbEguv/BGqr/J6Uu
mth+oD4CJayFIH7GiDlU4XEILa8gJqqTKwDTHaGiEzPuRPBYvPEFts23r9viA2iqQ9E570cRbqpP
SyxwY+HSpCN9bJUMUCmdwxm3jMwounBrbNx8ncuGrIKagNFb/PH0TZKYxC7zZR1IrQFTxIF7bUO8
P/52CkJgf8PiViU2uwXS+qCiDx4ZVLvEco1hSyuiji2EqjUYJIkBuSlmoZm4upUER5zG2rqqLvNh
mhuATIKZqnMpcROCLKbRKm3F74AbJCphbBsm/CZalJnr2T6UbKBZBvB0W3SVvy//ej63cN07k+Bl
4JS3ZZM4EkKeuusLOEua9eNqUdKNJn0vLvg7FgMARY1CuVQTn+kjP47f0I8roZ4r5KDgWInvGWqi
KiXZzAhrMBjTr6ba2MXMD2MB8HGKeFOrYqh+dMcucwXYYpMBpLlUc58uIykG7QqPtPKUZRhk7IpT
oV8cT+aHb31CEqhb/TFOu9zGDyFdmTLCYM9x4yT5CykwBixRrLA2cRzwwCrbEB1TdCMsuVh9JfYr
nZq7UWWe00fJI5rzDu0ZK1lE/c8tIupzTS3NkU7XcX2uRYIqSTAYGPBeQ8S1XHskozcAadyje9Am
MuSxtqREBCBTx3+r9OkROASMBTiJjrcOZdGsYTrkhYi0I6GbAUZt9xFqii09TwhvkFKG45pwfOVv
8jXppWUl/xUvnu9AzNVmjv8ERGfIEFiHksYH8HbnGKNFmXfLkkgm8rRIQuH9kEm+C8eiqNpJpgc2
b9WVI+JTtFmIaue0EQbIJYrmGhixF9gaE4KktJEdqiy8gfMiNcAURc9G/9zf4rF0JwUeLUZqsabu
Jl0wP+NRUA0PEWaSb6MtJaSzovXFzEb7fufbfe98o5RNtaID/gZpzNnQN8trd/erSN0nOY96zL9/
YYYLwuPsfPszp63+almArA8tK4Jw3n/b4yW7PuvRabz313ikWmMeGJwkO49S7nJhGXiICSvV4INr
G+ntbZwJleCrWe/FIItfMtTrkfheQsjmdBYmh6uveUj8IQKTsc/pMg1I/eb/dfbPZp4e2eWPy47w
67EhSOdmt2HkRq2AxJG+UP4eWHrdTHCi3xSkvjH4g6kw62e1654IT3AsntSxftxBVhQvvlSUmTHr
IAtkFjdWNSXMRNJoACKIZiq73USN+uhuBbon9fPiGlYChoC5aOoOVfEmxH21RbMGYSUYZDiOdYlw
Jq8HhVtVudVMhYX2z+fnARb0x1WUT3oACCXPSUd5PatBcwnDefLK0WYH40gD4hkEW41YzJD/R3Wt
lkLyH8bqS25fXSZ2mVSqJx4wnrwZfZhuua2yWZEks9R51sl3xadF5myeLoAop4WSL2C9Vbu5BPbv
5VRDiyEnMQv0PoH+j52FhJZEMgugBMgb6dztBvKf+X2VAUC/FT9QhZwGov18PaJO03L+748HPRMa
twb/c19bPYaVsd0SFOpGgUWj41ZxTM5UUjxhzBWMGETjPV/BqP32e1g3L330kWI4u5R6HG3DZRR7
5NpNkYcrmRV30x6e4Bg0Egy5lUkteDIwx/JelIxZOX60niQ9Si0hyMwxIoWrSPjy2P4xp2aw1GZ3
OfXm6KR9SdUg5LHdP2YebWWqwcDtDxjmc7lH4YOvoQjmEwmVz0EnBPEydziaUvtVwrfV1JP6f/jv
EEnzj4kPWkOpuFYIq9Ok6H+wPRQUVESC02e7UQHSZGB8BHB22odRdcgfgudlZizrgHcstdSd3QDQ
5qNbsi72SLz9ES41/LsNCGyK4u5XVEVN5VwJG95VEa3cShdwmgwRi420VHlAsjV/VPKW96KUWu4r
GNfaa9vQvuPR3QTUDdq1hTQlNpYDxaj0L1GyA/7ExeCR3qMfCbgDp1aT1IXUY2YPkNUrrd9SCwKS
N738nbV/Jk7tZEU2fWlGWi41klbtCxbM0QCNJfzY3B0+hZLhLTAa/hPiniTNNmXnxLNm3UtZmfpA
hn7QMaSRiu7kezNLTBTH6GZ5sCNTqhB6FTIgATod+LRvKPTqP8v2mR1RhWQW3GuwwK0ZRaNPjaLz
9gkvk3XbnRnEjjE8+H/P7/ISrPlOgI1EFSrTfxJyBICWdFxUzrUUzUNcpuq4KQC5fFvn3KHsKGhV
kKUFopWVUm9l8o/hTnoqwlOLOXq4aZ1BlMaFxpetktWV1vyOjZplGb+KbiV0GL5fcAsbV9D7ReK8
4ea+YP2MI3NVIazid5zSchYm+wCauLTqGjhOYQ7TCV3G/gCsgkWeYK3EA72v2yE8JRQqMEgw4aVc
Tu2B6klVcB78fRh41cF5ofJwC0DYnvHhlySrg6llR6VpjDxAK5zMeFmxeFxrnEPzNLkbtc6m94vP
nD5/KByQE4jXc8/gdHBpszLAse90E28E5OLm9XW7tEQsg/A2ppnmn2ci19Eu8PZROCNPjsy1wkI/
2Q37VK7Xnd68DUExuqXq/cKO0dQrsjjju9RflV/0pAu52pAtU3Xe4w7H5W6asaY2SR3WyGrVQ6dA
iBEVlZw2qMcoIkcDxIaRwBM1xnLTBba0YB8tBCg0PS+4Jn4/kVrEMc0YEcegke4ymj7lszySowlW
4RecXyAoNa3By/xRSYfy/2wSEEz8KIcmCDGwhxltD3TlrLkM989LqZQ1Y7XBDw1v+HuQC/hR5z/i
3twnd1pss/DlNZcKVHICRJMyrWq6AGEbiluxMu+0f80cKnSk600yyw9zfZy4QjnYwNwWKDvtG77o
1Z86QU7j9YvKT6G5HKc+tu/YL4EQez9b0D3LXXbEvSDIHHTgxUlvVdTc3xgLY9ob6QyC9bzWC3gN
7uj9ySsyfatc24mPdc3vwuNDQ4LdNfcGNKiGh5hEeBgS4a7E2GMOB41HeWlSHKkqin0A3jvC5WgH
6lbt8wR1JX2dBBa/ShfkY7pgE783iR/jkf2b9BiOLPaQZoCVyIGNrGbQyfXSaR7lWlZdwfMOlOR1
yyi/4a/+X4MjJfKH13KzEtAxioSpmZYyecGWDd/raSVi5enxDPEhy7Vx07Vxtj9A/qV0AgmDJi9a
XkFtiGwZCit83/e8VybIEhIvFWcRrSXd0OB9IT5ne2kxxPYy8mRzeTpU2oxLVJ8JptBpZM+JrLYK
EZySR5oFJOckm/5AzB7uNy+k/O/IzzKTbCsVciR3TMh/ohzh94V5kbV3lpQqU4e8Xdo1crByI2gQ
C5nOWNudylEjSrWLGCmlFUOqHsp403lRoUp08gxiHNa0MIwaNUoqmm4h8v65jOuQW0xlgPTyg3oF
BgPDgianzozCPqO7E8m2r9HvNioosZax5ESW7mG7wxY/xoKlP461AhrrEFuA1Ca7CnVkhrpruK9P
8xT4k29HXN/rDXoP9jy6IjkPFRgU9acwWfTBu2VQphyb5hEmuJruSvwPoq6mHPkfOgFIadtyOent
nOCkKpU79wUrg98trD/Rs8PBGH4u/mT8geMdINhh7KqCGmM316F4Do2NhAA7GvBhlcos1TtTmi8P
lHeZP+AkXApoDXAAvBWPubo01xyJQM73jlDy78z/76tvV1T5lA2cH+kustMQQc0gE+/EJksouK/r
QxtCpDbzARGX/7F1oINiroy92PejQi8KikYoarFiYaJ2rggS6HzjMmW1sqrSSVgnRnVns0hZcluJ
5da4CbqPWeahYYZuvZodj4sN0VFobC+UvdyqhKhyralFT3ZYjsjdlxZyBTrXy1lSnt2pCyKoB83s
6TTe3nVw8RcEP3dqX1FC3ooMCyLIaP/WdTM49tGaNfaF3Pkt+4hLdv1Zhxg+UsjYshIFsuyMeww5
l3U469f5UVsE3N6X3XchPF0hFxJnLyJdN5VzwEV5o1FwIkA+H9UyFqV4PIaeAfk7HG5bWu//2D85
4Uwvp45kgfRId6u5sI4Nqq6JDKVfVhx6VQqmUhzVga2unfEia/VX+DOY59ZLRAQ6BoXF6Zpfq6jc
Ihiz5dPZ/ABdXJC/Lo2lL5JIhKMsA1IKL0QoY7vkoK3obSGHLFIz98TKR+whUaLXRgdIcfKAUh+/
As8NRHD5FnVTqgb94/DkLGfCKhEWCYX1pZOtCK/Ak9Xg//OqxB0gXpbyz8VRfQZsry0U515eePuF
Xd4LOq6pnOQGwUqSuWtIdrIGCGnEzWNBbJp99ngfkmMAaA8fwAP6YkC/tHWv2alzF7WtyR3KnfM0
e/q2Pts8+fVFTHuFNUoYeAm0y5OUTdymlTQwfy7GT5REWjAzWRidNlu0gG887QZiNAhwnOc/O629
SXV1hRdpN9zRggYXN+cCw86p1M9UvjghTHuyGMgUJFwAyQI3TAV2Jp5/kHJurcZfKTEcKD9rYtEl
Ww/XUrvVV5MeyOCAnTbinGYvHxhWSeApmEJwnpts/XcfTOCQI10LpeAP8vY7rZP//m63YjgG108Y
Q4ZbhdDzmTAdRjwNKlCbyFKn2lLfeoVlouaI8Qd30y4WVsljAqGviSAC7/4ZcnQ2mMqdUJuNfBdT
zP9IUnIBphNWWLHBu69ahj45ixJpcBLfXdfR8S1TfeDusTCOxbzdr5KVQ4fIq+hn4h68lONs+Xwv
LuV2WMaVHMHW4CMMr534bLBtzp4IFfRbcEfaJa6pwqjseLwNuHDyZRCbnDsDVWGYoJnKs+YRhsn3
9rT8YV26msoDuIj/Ly9LI4H4oMd8c3MGE939d2AGnKiMmvuME45WDI5+otETKADdygoBLM2A1vv9
kW/7Kh9CLQQh/mnPUAAwcjtIr5Ythff/Hq4ZuuyRkWB3EMXvaQRLMz+E6k/0IXllf4jL6X5iZM3f
jKGnSLQNTP0LTCDAKb8cb26Wu4Rmu2jXANr/vLjJhedlcSUTSzqwEDEKSUr0NkqSyMrWjxKVBzX7
KBcTX79bh7I2eVRMMSMJ/GEgXDnvMC+Dspw0Iv8ln37fXetJH1DVZtgBYmv3QGHbbhq2H+vdTnXn
GGmpyehruMUMSLWfEh7bmE/jKVo1qfgsFwEvu8mKS8LqkUWA2lr8rZZU5ksin7bSKRGH1JqVv+V1
IsRse3XOctyMDG9EilDVdY5uDoKCJaHY7+LkqpsUWkvYHtqpCUx987Zs3I0hWy4Pb6htOG+YgSu4
2EcXAPBo2VbbUCl55vjCCvfPEba+1jSF7W/Evxqa8cAuEpyzSuzQCg8cH66tkYaD/nCUSVObhDue
dXnYbrUHC6M5AZVPntpPExdChjqi3ct7Ywq4bUBiZkWkr8n8hhsoUWsWGdUJldvKHY8Z1sFrvASF
0rtGhoRuMN+ogN8FnjJiPMmgOYp3pzHrDEW58r2SDHZfu7jOtR+vhcft/NnvIfO+xMC8F6qZV/xb
vw34jaxyD7stgRuj/gu18DkJnlHdNxqnj6erkRN4qrLxrPIOaRLINYL1o5bLvkV5D5qUiwi/X3hI
Dgfquaike2HM7Nlti03BIfPlFTlKVx9k1n0CmdM6SsrLOysloccnB6Ly0Ljcbv9d03gRxKzBHB3b
hlKS5Re45Fwif9p19wfGuQeY9C4qczCvtJg9Kqk3YZgMSTfwcy6Ut3CHPzZihHEJUpH0s5rHsvGS
F2AdM9aZG7l1xS4+FyYxInRZDAhzQ52YVifGVUqaifxCnh34rS46ZcLc487VsdOWeuPTyQANLDQ+
yA5Z/EzdENwg7K81s7Ur3kgpL4HMdQRoY4LnDLH+eEL03evskBOE2dzrdSneBLWESBXZExZCLhZ5
QfFYRTuYitsH3RMyvWJvIhQXjDB2Xg1C2w/PYDo40BW8xZAcEmLZPe8eTOgUlhyWoRZzX3pUGZpG
YcnyIco+VmOAu9PoCwzUIWCfZ6p9FT4g71wWxrp4W3Dgj5kJx1sQtgWsfazM4rqLU5E/oD+5kA82
dcnzB9d+fZXwxEbzGzSTA92npikjsirpowSeI7UjH1V4oPX/MYmFYxy5a2YtKseujtylVNGmKNgU
tHKwQJ/L1G8K8LclM6yVuBLeE0PytBFiBUk8agVgqG6ElA9R/9TN0nJYX/RW5ql+olVO/xY9MKI4
cPbdEYRwv2epb8g9T7l2JYI9BE+qO9vgNDHu4mBZcpf6DFNoWB2TplSfzkRGFxva7hHe9nmLaGvZ
QAuDxD8iPkuPv0zYlW6MtC4W9/AauD3Vx0MfEBkZjhy2gINBYUE/hK8hKqc97hp4uTQbPrrbhkdT
nq60hTPGLyF+f0Sn+OSeHRdwfywnL2qZ/7n1HXIw0LO5Cc+BtospovuiknvxExMvuhdt1eyDloDp
f2PdqU4mGbKBsEpqyVvV6UaDtAH03GuE57Ufb7Xi0gmFLwvWAlXNiIkxVc37pL6pkSNTGJxhKQ1q
fwu8wanjLjexBSpAvl4k52l1wYcZ3avt4LGsjADLEKMhRoT6dVG70vYkg2PStkBkKPuPra/Eosix
yPzH0FlVM5Pk7Nqrdy2UzJxdSRa82iTegBaDOHu7bNUIhuz+UKDZ7/bKGQ+KWslWGA4OL1Pxkxzq
fKeLNfDFq7D7B4wRJnSqfCFj/xEZeC/eJq0mfnnRDWeCr30O+rK5PJZ/6f+S1OTck6svyQIaJqQz
ucpuz3cjP9HISzmI+Bu/ceCmf1NHR4lQ8xFvU48VndTkxLVYwolxSmxNf23OlbWYXaE7/KXoO8iF
XTPkXhoRQ5mO3ILFerI9z71+z7BFPvv2aq/N7SubILhZe5miyx7N2FBOEWMV37P1CDVJOOelYUZb
b48kfaytALByyk17tqkSwm2mSe3Zap3YsWhilKnaYHBj3NaXgw2/AfCMN0wQ2orpQfNfn0GcDnIn
B8cFkzeumwQVK93B5a9bGON8VDo4fZZZIvVHby1lXiV93rDAF877HJO9WvhpOA24PvrP4xiaymzq
5OKjAkzS43AZJFdFb54tSsW93DCWRXYwDNcRHM98rr7Z9sgDV8vH/DL9C6LWEQ03t43hKzlinorI
HBb3mDCMA0CJK2IchQH5MpdZfztp3CVTTn1bHDF3/3WAh0Rm5nwd0VBrdxE52W4B/5ybHf5QR6T7
SiHmiwnxYvioskJwShAveR1L3h0Ggjdz6sQ9Zsz9iyvPrSLJG/nXwxIhd5p+nEOwLoEY11NQzJ33
fXgj6yIoJksJ6ouSi6lPufpqknfV7Q9S64RViBs6cU9UekvUGtvJJx6aMjAguRvqlaaRrgPTw3/o
0xEazRigsKg2tH6uZYw8yisSlb8aNOF+mEWrvBJCW2FK4zOBhrtM8YR9jhHIOKFPFhZcvlOAzfTs
pG+O1m+5uoQdEsd7KZiwrWgLueshlpRq5qHta0SxGGN3zmb8tlFmcdaW4UjY5Q0Hqs6QiA42Wldk
e96BtQqNXh+e7kjLYxL0KCXD5YwFYfhNcwHUzr3g93wTLb/Lef6xzhHOvRaA7nD9lawfV90fufV0
807rxvkCtHJidENxLeYRgtcZK8rdiARxHD/4hoVcwW6qSUUt5sqBiJnrGwttSMZzC+1WFqBCOy/c
jPsRSEYVbn9WP1OzzjjQB2delGMtlHPfX0TYUDklHFpByQxRQEUlv+Bv+dfy+itlusq6c9w+00DH
ySRZe9jyldbvcQwKVCcp23USQWBl5Fcctr9t/OpnjIEOFMCUrmuUdV5YMe3dtDDNt2Z5I147plAY
/SMmazq9Kl7SNIT57mXp9vDav6KHY0szZ8mzGM5P2bzvzOkfcrzSjd99p4nJQXh8zA8cIvaG/s7D
Rndg9Xs+QdNiFcJA65SL/9dW6b9tEp/dFbq8tlKwkkcIFrFsJYp0QDZ4RHXBCkQw/W/6bU7Ly3hz
x5nZYt0hNXcrTY6x8/BeRL6fy4SKFgpSyHUoiqH6zYT5n6FoO4THAfHCN5TEb+S+FUO5iZBJOtHE
354+UD4REDyCz9DxxHTYUkq2TPpkyggIWfixEjRoetuar+jT32sYVIIZZhQTS9AMweQrXS5kHNW8
VimE7IIphqDer6sXaniG93bC+ncH08lQ+kzWM7N7dy1DbG+v17iXXkZXMzW0iOJ4znPxJXKhvyGK
pYAva4uK/tFM34PvcyJfNI7ft7NntON5Fce6qaiLGkm9HV2Nn/AkxxmT7a6iyNFQlfEegjVoJxja
dy5ZcSn4OwmaLR8fa5a69vYAFbMknSlCvzrjymZQjcPeCZAvVD4RiDA7sGvif3tua4MwGRIxJN84
Qb4X6YYZnFa9sxi5EVMr2UoWPPeUZNMPz24QJFoirBRgi5INK8WfeO2IdCV90r6GM3Vkmg1Heq7z
WgfUeoIYZrZhFDb/w6neyfyeoKvVXV5oV1MyRqf1YpEUBHBryUl3B26pAVv1hf5CZZMEi4/rXvcX
aMTwXudun3li0H4ERsoQR5aQRd5MBIcQMLURKsNPdzAxOXKVPv8LZGlo0/i0yw75BDB3VQqTG4Ph
WogGN+w5BqEDLZhrPXk0VwfG6Xou2p8sMOfx/I7lkRl9IzcnAP80SlvhYTQUNpAK02V4MJAH+1nN
YJ5V4wFNuf6AUszTE83J5azGd0ADcZn+ukbtGtXjIx02Ibc6HNV+1+uEiDaaPKMO3AIjyFGS4FtG
jblDo86GZe0/3EHXKKIFunr7Aqohcy2YmA8N8jRQ7ACV3nMRH6kpoQ7kinogMg4eTAzlSOqouOzM
Bf/kM7Vx1CbcHquJ6S9iV8YdT1eQG8aS00IKSSXGaivGLPgbGMLxDCehaGMMGTzPR4qaWXu9iDYW
8p7fwmkPFvUS1+MaFw77eCw9qso4v0rW73t6F6kH82bdNUhGGLJ3k7k61E3UM/gWwNtv8fNdvSEa
dB/3/JpXFk4H1TagnO5N6bArydDCLRhW6aACNNPS8ANUEsoAgP74f8k7iQfMZW0wOyzvK3zumus8
IblmuvRsC+qd89rAs9c838otFyATTvkQObhwUjZq77e8hlG0HIxOQ5EF8dEg1JaW58BrOLVnR3ZK
mNNwKnTOvCRk0dkPenXyzsCGd3a/9dBVGQjlrNqqRTTZTRNridZPZxnDbFz5MkQyxMClpak9XNIJ
8OZIUs1otpNG3wYgJLLPmrsL38vrt2N0P8muiyDf3+4NYp0rZpWTGbTOA4twxn+Z2MEyxBDiG1z0
iuFL6HNslC7UJfdVVIsVj66rCHIQRNOCbBBLlkq5I5aayv4hB+bNVoHpTptnFrENfJxiuP7OoP3m
o5CrUI7afb9uEhMspu61bp5oVVwYTeU6bAQFWuQqJZ8WfD5PVRknSQuby4EblarvRHFUUoPpkDWN
Ri07xnhiLIWbsKSxFi/kts/3fXjJpmPiehZt99tvGnKHqW24k1Qr5RAVEaJ2idHb5Yf+ZnS956NI
u+L2N2drPQZYL0loKuTN4cv0TFie1wLoakUboofOZZAFn6J/EF8CZBkapYeDfjcmwkdKwfYYcIFZ
B1mJyg/Bosaw568K/WFdpQHQQLXFxlJhnJ1neQCPLgKmTpIcH0xUO+NMqRFkJSwVXmFvnWFSbULx
NYc+GGPaXj6qJkrb3BIEpDrnIkuu3pvaM1qVihK3Gk40Dvxgt4rLWKAyFfF5PDzkPSzW6wSGQbAd
MtbVjfV+1yN18J+36dzBwQVKCW36/XHZPIKOhlEXZ9TM1/Ce6HHYd5Y/0AfpNkr+EzB9OauPL+xn
xnB33Aunq/OFisRHmmlfOCFwZbo8DSnxwUaoGnCRkypypCIo01qcUbz1yFz2k1TQfoYmdWsH0Kda
O11fQ8k3rNTJtBvi/R9tbuofqvSO1fqauUqTGHCiuvPFbSi/N0FQ63f/2WZJzqu5tct7fyzwKHLQ
QdmAxnieC0h26kEPYkQlbtc1PkARQJL0ZF2CBqwhdeu4dZQ6c5+nbBe5mVVLy+kuguzwxC2rIOCD
sQ3nUDxTmQ9oVIvz9ZpxnWYNDdtg18zIuF6WlwbrIOJPUjO8zDzE+vCBTPyH5ZpBWlbSI8uSAkhc
3e0As3AGPli6x+nY4YP0+Kb2HSivsgSM6Ad11H3nv5UdxKeeORjqWucFok5kCDuUSfvH2OOUKBGs
RqLUTKupGMI2elkKWs78K23nkHkCmEGZOJh9WZLrWZ028ojph0rXvgsbi+/wCVNK9FvOZ3nYfuAn
h1a5i8YTzmcBu8bCgFDJpME0OVUotlv5ZQyF+jET1T9Y1rqRkckmc2TZ1SDN4xkjpP+0GVakU2ed
BZXhq7Fd53QL60na3BgP/Mz6Y+hpXaE07QCKh26ot/+To4iDidBX0imuEtBw6b9NHOR+s16EUtKH
QNFaHfCNIAHNYf5GqLz8BLHNUPKVHr6MEFp9ErF0xHUpHRdLkTnvYfciCKwXz/chi4HXybvXChXn
ouaeu/SgldLOgpE+3kdffI1V8CH26LT05esQtAgwN0WuBsnJp3xZV3fyfWIgmQaTruKNxyUPyFo3
vxCmJgyJ3A9kvTyuBc/TjXaFDeqr6ZOMvYzXGKmBKpP30sYGHE7xjb+p2QxhPnKx4WGYP59zJC1J
4Xyqe5mCzopsFCzalvTpi2IYYxUnZLP/buzcbfcAdpPqYoFIPDYwExvaiC7VMLf9gTwY48AMQQ6C
vWjWGYoFVKt+C7W9LHfHJLYSVlkHwmGDoPvzw0mILLCKtKfXqyaCe1ZbOTlKWdU87djkiN3JdXA1
fy+W7Ofm56Z3sWpS0crtuPGVe7ONgyQz2IBEQaXtI2oUbyA+ylff0ufbYCcNwvzNKAJFHPClIiv9
n/KXpKZHsKHF7S0N7QXpx5FPYAPLBYSEt70taxGfpdLgRxG3yPCHMEjURkdvwajM1BJMSlXmfvsV
gKo79LbjTjbaa+jsGgL4OXtc5dfy8wQNqoIcVh8V3KKyelRLSecJ5ozVPqI/ServC8z6eJsB+0Ke
ehRP/mmi6kKw+DwhK4GdEGKQlOe9fFsemCHkyja2jP7WkK2iQC+UaCZKS9shmCCJRs1Oq8HQiszF
sluJVuQjFPrJ8hMkwfVjzrKkhYcLi24U42DX++0/Wa5BHzNhG4MTwqfOV8LIhHSU6fN30t5OlW/e
tIlAjPk6fEU8aQdGVypjZCHZyhTF5l1O1sdlpFHH7ui++Y4sQGL1auQ6UJQx8ylknqGtEj/p3Dmw
Kb2YvhBgX7vjr8ZSGB+YYXBwc4Qj7Vs67PZgTzxQj1xo+lJJPcUWo+gdCVwlYqpYtyaaBRKBYnXh
j5ANhvwacgt1LVByt5UsgweEX++5UDM2WKXD3eQAG3dsy5mZWGgNmQ9cx4LoE6lKtEwYKaNP2SLP
z1JRNioPiLJdP6SkeRuP4RSsvTDWrqtitVurWxoChA1mLcyk5MgW9SsVxn74QFBQMO3aTalj9x82
IOzs2L+77EtC/0czSlz4Va4aus4u98F2d89ffDYtVt/LLgp5YKgk9lpL2H4Vxy5J0+1NIT90vYpl
AsY5qxLqPMpRYDnHXpg10+jXjaUylRCbpUKdqigkVpvqDLR869oAY3QoOQ/9A5cIN3TFc3d83S/I
Bb4z1aryqULWVJNhPEUNYRh29JsHlomOkHuzek8x39YKrRy1lWsIxT78K5NVf094V+VEy9adm6yB
nKTQLLTevEnR+zNz9wfin8XJYFHlB7+TinoIpvMfUZajzuM15GlBxjdalz89ErPbb/WLV/6tfAiA
AtmT/8uBbLJSbxouSQZspLuw/GfjFyfH8uTzr4usQAG15rYPqsg/pbFFD1EmjVmFqHLplaOJM71T
5GepeVM5dBh1kaTviRRA6vGtC897z1nQj5ryvJk5xPleoQkCkRbs9F1M3sGifUQ1qjuICGF01zGt
Gq3tPP3BDaIvvnyb/Hix2UZLLIbYUK5gD6//p45RRXcnvNdwhEDb3A2I5Y5ZJNkwUAt52lvbjeiF
LnOQVxiXQQpKbr3/c0iACvGzEmKXNhOFb2MwjU1DaJZbyalDZ5299oSGWtqeY92UbFgfvGcMLMxx
H2+sWAZmEJdK/743SZ2uTpJk59IrjiuT2wUKndz743pSIIwsJpsLRGeYmT1arSCdieBh5cHn2/1F
tcKPxnBaAJ92fh1IZI+vqWELWcvt+GepnawLHqVgzNFADdk7CUAGEQt/nlY0vWFl9oSFQ2E4xl9n
iJ9HsyKYrmpLH/1taNAPJ4uerLNQniAu6vbM6y3VpPN+9RdySysLUiQmbEvRFtTDPfHXl0tL4cD0
uP06JK7sIoSRD2Vc5ovriMmaqWVA098ZDdGeRfsFFCSZEdR3sMCUWlyMHHYLOwwPVNzeBXTJ02Ea
dyBQGCIFy3Yj4FFlvj1u6mMjUCpuAMJIMx6SjTjp6s0sjeR9prfEaS1os1xKq7qS/BAMZIR3KWE2
cLD3JUYcB54tQc6ARvTYqz0dNy9KksSxSGJc/9VZrLTFRUCcws8+qfa8z2l8SwuBNmyiwAF1QXSV
nW0xC+4daYsQAmhX0UxIhpZztFY0rfDeAwjarbwc06jwqA4aS/x/+I0cnc4Mwl/n4x2Qd0XtmxsN
LYmGLdve+BPWGOq0Fe5N/DOt44Kr20YxD8q5SiKKYKlXWfw4D//T7qjiyn0ObUHHvYm2R9Dx9ykE
jmk4PLfF1LeoBp0RcQwKin8f6DxlEbwBLG2dAdl9oxGLzI+zRnfQfbLcpkWXZsS5dB3xDeVAtvb4
PrbfYvhaxbGnec7llRwigD75bkc8bLkpfJt0bfA7Cu7RM2/G2NI2oEWordfQqc/cmXpGjqt+ArL1
Nid0E5gIno2SopmTb4ITmn9dTa09UEIx3QhKMM83Xz4Fg8GmUsRGVFfIeNbLscjiCMN0oCkEl5tA
dFWU2lWEplGKYd+TVx0HjN7V3kb4si6w5AlP1246KHkCxLZ81Cx9QAQXMcz2/Xo7OhfE3w0HJOAR
Uw50GZgHRp7qvr9vwATxbpKr+KnV5ib0MDhiPic4K25IbJNUu/Ex8s4aQkJcXKzOaXR/8K2L5eCS
hFlTkZL1MN2Sl8Zgn5u4IUR1yR/LuWoPyUEeB4zb9mYheqyVCz1ZGCO1deQP6+EEH4oqatSfHnq2
tuDndwpZ6Fy5LB4d+8cP4+8SGOH9X71KY6dbbwphZAdu5B0SPcWQn3/r2ie8s8zTJiJ/uuNkAW3P
7z2YjQx5GtsF7W23PjEoQg6Od5EiJiMxJrfrnqqMsIyd5BVkXhQXKJ6hzLsxinmg1TGPipl/06Wc
WdaY6PnmT24VxCbxxxUn5wl+EmP0cf7jMzgqSPLtGjl34nkKky/Syf0vTQGCjG4+5vV01BTDoWUh
NJQUrhtRtAGGIAolLt7z43AEeHF7vv8tSblfC3FOtwg8pJz1NPKppgJburAEA7h1Y0Jmo8qnBfWR
ZDJH31YiGh8hAOXvDSiH+QExwj3nJMO6ra8HgCGwrFF0kaRB5gXF/3iVQ1nnkZkxbuM+QnPQw4jQ
6xvsyI2Zn8DIQa+GPhQdoRrCQBD14uwgdyBrD7Usxz+Sj+K8btzUgRFCDJG8Dc1PV+xgmazF+Zvz
9I687jmjqPmMRDwBkpUTzlUs40m6FyBdADtSoZcJR1FOO580m9MSXPB7PR0RaUoRB5KZ2Cc+gRke
eq04h7KG6xgqLlWREi7Q8ZpvzSxQDTic2PTnaXpxwUx5QOUL7T0xw06JbAgcFOaHmaWlBbP7D+M+
wAXFruBW7RzoDN4GnvuPC8NVT9YTipb43LZnksJDsafA95xB52+cXEn/0m9eUYuRyHe+mXOPvYyH
2meYknxQGsE5G1izrc74qlIcramg4md42gw8R7lDMZt4+mfGaD9N7Xb+CpPn3uBscxXZGhj7QcLn
n8Wt7vcXWXFF3ojQJVKNhd+dY0wPCqJe6G0EKzoVxa76+e1CM6AUhBOCE8FiKt3U+9PqC12evT2+
fwBy+7jkoponepm5YajrLVzfhXu+RTwtinfZvLsnND6a888ToDWaafOhDSROh0qHHMYIfgAaNhmG
JtEA55Gh8szK2TJgREef+ITeQTQxZpcBGxqBz4h8WQVaBZ4P6OC9KmvyHy2xE8OUvtxjsH5eli+j
Q9vFNsyeH66/OdDCfpDzRHdvooUMbqz6PU/VvIqxEIDayI60C9B0WT17GqIQ0NyncudYE4Oo3TaZ
E8FT2vf/2JZENQmJyy0KKNfxCdFGhpz3SqiWXzTb0cR4+69BFVLG0uA0WXfZh+vw62TMZoUo7B0b
5OnLLdgxZ3ORwWa5O3sr3PyDkWS0kEQpceK1P4DpTEejKxIWjGV0f1jzkwNhCJ3PZ1vJd8wPyRJ/
gRf7se9DhCmnHhRxI4MZFCnKy+uCZJm2uX3jKJ/1ozxuRYzpvUZpvwo7vrmrWuGcx/2jzaaL50gj
EegXUSpAg0SGv23z34LwST13D0jx3em5WHZ0amn0bDhEVZYhSG4Am3jmiOiW234ggg4WwlNO7QeN
zfrzsP46P5ql7Fb1MoH4vJ9NqG3i48jHhGFbI0RRHCIWbb5GjalKk4naSuNFsmmqDzgzg9DzYa+J
EwxwhHtZ4DdMpZrwv6gqk4p36nfmLSDhbWEXh/u4RQgQzdJY3Q1+/cvSiyh71mSEWhYgC/yItQWS
ku0bGTBx+M/3D0JJsDySPzBtO55oL5o8W216mizQFV+/U3XsE7PCsvrl1XZVBda/JpYXPiC/gt3w
HIdFALLVX3SoeyOP70UaHESWAWwotwqrcocq4274lu3CLvtUskiyb7fjXn6S8TshO1p5aPGSJU9k
mys0d0uSGYbzkDZ5Pe2FIJecMWAh96iiXJOIW79MwA6Fe+XoVz4BJaKfeE0gyjn5V9icDC3+LjZw
5D3D0MOfYlu7LcYgcpTv+BYPTGplmawo1/F0uPY/NI9uVD0Ddy9r/4SRKtW+0FTjXcOCHhkSWtxX
DpAXYN2ZP4CgpUVa/k7Sg4wjmknD43lE6RXTixFbLgH9MmXQeMD/llYqgYKBW9ueFEkqBQCHltAe
+AqRBvUlcNNDzTxsYakkXc46ZlkR8NGP58G+M6fTS+U/AtaAXW5ewYIP3wDtqJ+r4cMe9SmflJYJ
i7YmtkwjaD8Jy+89SB7yp+03rE2vVVjQotuOl0dxgHi+v5c6xQUSvsfyqYVHD3dvbX49XRVL5fe2
XZh1KL2O4UtmgIzf7vDmYRU+wT617ne8CmQo8eB3ateyqHp/vVsEZlNuNWLFgz8wEgedRAZP42Uz
9reVru/hCmleGJOavgfUzx20SBMYucypgUj0KPWIl7ukUduBW0f4DxR3U75bUatbUaJky2FzJpzz
3SmV6XQs486OfVvHLUXfBoWfrSQBXK+hopg4s4hUm1mFDR42g7t1zx+oF5X2j7TIM4GUvx3YPxeZ
VCMKmtCR+9BsMofqn+tzV5UCqdiovcY6bgYxwn25Bh5V6+WVo54jEFP4EWNPaUmbZNmnrA+eSgJI
CroZB+ExUBY8aIynzTxZAgKqSKvmg1SyJXvkM9jPwosaodqDaQ0ESddP75H50vcmq4d2LtLx95O2
V93nBZaU4sssyXsaViJtyB9lb53kh5ZMd+yYPLtiVcPJ8ZPT9DZb5NctwvIR23lYxx9yD1qAeXFs
8DDtFQSOZeBAvmkuuXUDHLubl8Eqw22SjIJEMemfgU9Gs7Zxb5V8CCmQIUwHiE6PWIaJ/vqH3PvM
dYoOsod7ktdzDnkCHxLUyJdaNP8xVs4lJms3LZReZqgsVI2pIpvhqyWIZYuVk6Y2l/rjqJLY3dYo
UobCy2IDMQyFs6x19DXxllgqRapQfczabqNDRji3xpadcPaEORXhCJqEBHHsljH4Jea14R3rTVV3
L9J4sVFXqrJ1imvC/m0xD09N9Vf/jstjrcpwunGirGuJBrUTZ+yWE3JTSSV1UxxqbQn7uJmkV31k
a+CoYQJkB//2Nfztws43OiorrMqB4r5Cw7DNYMjE+Vc99gUxgeouHnzxvQzo9DsyzYW5WKXB9iQ1
BBK040v2gius0AKCkP88mvcJccy7kcmbuMjsrxDnzDkgvB1VevmLvXq+QcjzMDIV/2HnnGIlJJRk
CsdtWyytEABgCrxVzxBRkoDNQYnAzp6Z1pJJCG4sycpxMCdA4bsyJAj4fi2qzMYPpnnNeCnoUqVB
Zi3szg3mjAJlCDHOYqWoOWwxlFBBRyCKUd45+OS2UAM59McDQ5hEo1/nd5Rb0CdEdyMiUNPbkgPt
1VSD3xwbGGKQbm65o4Bn9oaOvh5oHUzgJLlDhWtPmUltAdhSOKDzBgzBA1uDcgIKdtLCMd7tTT6X
GSw9Kj7Ie4j5RmuFoQfVd1lNfnrxBxY+Ym75KpYsNEaOLs2JSwItQ8A6q5BENMRqX7tV6D3CC57W
N8gitaAyjn2i/Vd1reIA60nZlaGJXRTWZc177RqutmzwN5FCsZnr7wjKnFp/ek9F05R31enYipTl
XvQdbZRp3lsNF91wIR76FfmjjXBuQPRnQq0lG9MpWFZ9GaQFFb7Z1jcKvUlwc8bIOFilDZBnRl6V
jRiG0SIxO2LugC/yls+XCDBgF4QcYL/0VUxA7PmrHnjz8eTt9Q7uRHcNVDqYYuEKNux0qf/oNQ/6
3ZTLXwm2DnlnIj7DGtm8GdvJEYxTKRlxe7yGF3Iv5xbGUKVXdksN9lsj88PWDZ99SRjKBDoYM6fV
dsKkfegMFrWXmg3h1K+6Ubjy8jouL1vGxkf8bYJiUFqDkwXkgpPZzryP2sn4vyc23hg5MPkaZoSF
7R5W4hxTc7HEueELAgddz8scNIHxYDIjluU4/CxMJZ+u+OKAHhqqkUevMgjUx6Wy6uI+q4Iv7uig
dYenJFW5OWNZhBF++/ug2o3ogutpagw28uTL0zC9Vl+0MlXuSi8D2Xgi4eYYGWOWAqbKYW4bQfrA
/tlrqXCSvpld0buzsP5tFoVC5meV5ILVsmxuzTM5h7yPiYFgK2ZN8hVDU8Zoz9q0X51rZpicpVyj
aKBX8wIqgi1QwQ73GWBuVR4/Izntm2SQoj+uBjVWgEqPbDEYfkM9j2uZ5aTcsHOY3yPYqEJTB3WH
sTzCVZ67SEgz1eCh4zdHHjgOv3U0L+L7DQdDBL6fK2K68jeIwzXHL/nUlFwNctC0YrkKoELeZTZr
BMUcvmBPhzCZaQNlZDfnpU4v5QlYg0vo0xEkyR8KgmIWZdKkytosOeLDi22BOvrKni6DiYi9zTiE
Rs3XeC2i7soWtc03e9/RAF90oGsB8eXmki0alBbY0NclwH2vtIqWYLYzQ+diKAQndTq0LcoekpZq
9W01OrSjMN50ailKrgea852x2fbB5fbSI/SHf9aLgIRliynOJgLr6MFfehhQxKJqDSduqR39vgW0
4qN+8ylZuj4vDtZ7Qxhe34VddGqJiKlv2bVYCzhn3VpK5xy+2hod3BoGpMddLgtE+gPM3iMkgm7+
1k46Gyeqy2dtMT77Kbo6jFutUi5gLiOcD0X++wmCB1uuc9fiipLjGjiHqMaso9Hgnrh+DeCz9xjj
epd3qdYxhpgwB4loFk3Uw1L5iiJZwVFWfaIE8gG8SDfhwNi3xjSDD85/rfnkF+h/oFAx2wmIQeWv
Og7G8OfUFqNz1reVS36o8Mq2wNj3/vVwHTM+HDT7Xu2w3Vjs0lHTiDIm/6cWTWZBCyDOoNyNPdtB
Jtxdekaz/0J+vlHAMNBjhrovfn0oEdYpcYz0Fr3B5Cvhnzuo28wnUAfZfZCtDNSF+67Hys1e9JGF
mFDrsWkAoWPWOXtHfHNPKB2Ij/smIeFNWyLcwaZmjnvjvwl7ZnbqWva+GQfPcjsW9+9Q/wzzIBFW
DLs5jKRfbj83RcTbpbw0MraDRsjDJMmeo2jDk5Lc+Sknux7t00h8lO6cRvFKdQMHk3IINm/zdOkE
spP/BJkmXBg39mjVkne+hrYQu8RARiUI8fCHj4eLcRi0XF7AZqDIJ71H3kmPOVCWoqviI1YQDdFg
OKL9Dn5StYHxJvJvb4TZ4qOmAGclK687HtV38ubnmIP/CpAlto0O2BMHK3xSgMQ3STU9HsZvAWU4
lJ1bAAmtVrdziXqu7djIVS1fy37Gss9pFw8zehgGM0+FIabnaEMS9/324hky2qpjz66TQcvlA1TE
BBYqnmXtN2XjLqtgRM3URS0NsgkzW/I5xz1A3Z1YXPdk3GAPJC587EWj9z6WunXSacPNLJPE1l5z
+XggT+O9aTv38+NgVkpjOwWMxp0cuhI7ZNkx0zIlK1vSE/VrYVXSDay4slzUs9Qx4+bI/NQtHosb
rH4v3RBzC2Y4Pglz67dPYrZ04B2NpEuA80wcrs1ouwG33uqEzl6TZVdpYdAhgodU8mR2xgiFwOZa
GXq4Herp8kzhhVnDVZXUjjFo2U838RXAfi0iWGxUHixXwSHW8QzA4k+kLrsdzFCz7BY8rSYkTrIq
lYIUxWf4Zl55zU+dD4kzsV/V2E/f7rbCljAFg/uqp5LqFDvRBzcGSTM6QKrEnZiJ3ietQPdnfKC1
2ONjUiMmNEV/BQ0tz84KWattZ7hRqyUD7k5XIV+tx4RJb3ndxe8kD5Ou58KDS2vaOalLKOK08959
nTh2JWLRNG823tYFc8LTWmBleZJ7ERzipIGDR0HE43jOxvgMoVHWWbm7GfJHVCYQ3PDlaJd/IeEw
tCEiMAEnAMh36sUphYZQOEYEWX49W+fmTs0BYtdwsTB0p7C5UAki2xnhMxoRgtsVsIovnDrl0HCg
m60pQNeSITuBQvAL8yL3ATiBpAwRXJgVaZjGlec4yfgyRIV9lp3uIoQeH72nTbfHotGJaD6+liAA
+q0l829JL4DWd3rK5JNoG5S7toaaQPeOzmsyCgLn+yGFA0q7jM6uiMTdtbpYzxW/K2MQC57yAEeu
nH3ffRh+TIt8Ian+0MJG6YtijFs4QheOU6uHZ2vjtbNtS1+jYqXB6O5QjDrlOBgwo/oJN/kKWKe2
g6zxe7JS+KOE+2QS/72K3rfyyyJLrpqd28LW/sSnHcls5Ii8X/G0gMQMgBHtuLn6BiBpL87QOP3y
uGpBFne17YLHskEX3LSFrwG9Hu574wVOPpf4E/gVVuza283IWuHy6RdlDfRkDu7y4RdmriINti5M
ZrNfjYKO5N/9M+VmVNnJJkzi0I7BW3aLVH6FjtCZjx/cCYSiUhN3aUS/swrkP1BbeuwX/M6ZoEk8
m0VH8GtjViKb11+xMe1OJUeT+PdJMGYk1BAiLlFPSmngtW5rU8laV3UOZhm73kkHhU4tzkL5M7xK
DwVW6HS12uwosf5rvvudNv4CA4+6J17BPbTsfNpMaqJET7bneAzaQ10urP0fHgANvSU7zgpvQSR/
1kZrBJILhP46GXxW3ULoJ2YEJZAF7C2mYKjBGXAbn0fuHcjG9RTySEmkEjggASTV8pyaTIS0K/as
KTxkv+xX3weuertK3Q2w8QmiM4pVAw/SsbhcgSC20DrifVgAG7DWOO+TI2BXjEbgzOZE01b1AYRm
NzBYSgTNFY61P0VUWvzUxlBzxFQTcmmq6UlD3DtHXgOyU+mEJFHzgshrar7OWrTimgij/Yr8vG/2
l9/EromqbsLAdE+DP74HAcC03OHQUlBL18jj6ACoxIHlixb2JQCZVEx8Wx1JeZD4lnf+j+fE4YV7
CNc0cKFOVstkkwSICG66pQ2Fjx+mr1HzTl2VgCjPaMGsCaf3Ty+UdkCu3ct98jlcVxHfrU2RDaFI
ssy52T5m0igsIshnr5VzdiYQoYx9ahiltghfi6kHo43lcHEB3eUaB2ULU4hIzlml1eMjlG2vpmhL
d7Gf3dvyK5Yh5goQ+d1foD7UxOB4iXOhkwlnZ+ql9Y5xgkWC8d0Ge+YvN24pMAQB44yoKEWoiAOi
oNYGm5sVeOuDGRtH8RFn+BdUhpkdeqtpOOBooSCIvkpViZ/1lIu5sQLa3JO4aBO0Ba+6BwyZN6fm
ahAi0AH0Bk9kcwtQqlATA2nkNbhAj8zR1Gc57841OjbYA77NPiynENrsX6FsGOKO8M+SsDAp3MRH
eex4qgwQHjkxksNiBZNlLBkDtCz68OOFn8b7ZqAO4l99cl0sfLjY3eBzHMmNHOe0bEtTLU9KGa10
VLpt1u9XGoo42nG8AkHaCJgqjaGZtgZaGcuBb16vR6MiO1dqKxlcSBAiJwJIMcfo9tWZsCpu/ZUU
yJZwxqs2T+tqs+HyTUyVOr1C9jLOvSTmsWy0IQRQIq/pweMOTx+BkDfQmJY3y23sY6tg1KhfYipl
MXds1NJW4IarSFrjF7En2dWFC3LxM79v3dnO3jlsc0x5pk/CPqJ0/Hlr3XapKXCN6O74Pv1GwET/
jAv8DXmM7e6GWgQsM8Pp3/4KzwfLhJjw5IzEtmlPx9rinvASxO6okKRwdp8cwVvHsfSNF7xWzVmP
ezEY2Xm96Jc2A0AhT/EH1iRGKkSWra9ziGPGh1c9dMY6AFGiqyJW1krzeSSbMnGWhAb4X50/bvg+
QaKg1KfuShzreW49VRNhv5SA44VWH2D+vvJfZZN1ZO8nNRNFxP8HEeC1AaVeE6A3tbPF0faLZd/3
ZPwUJn26+HUFk5+E965yF7w0ookyEeMeq6A5loZfWulLIz9Nlv7G2IdEHl0scX1ekhLzAZWrPp3s
l7aZp264PlS1aC66Piw77rHNI30hZxFYtO6drL2jU0+e/oa6WVu+9Pwd658ltB5OhaC56TSmnck9
EXj1uYNUaIhrUDZn4flJwjExUXAHYioljuN3jKGPT0VlbrSBRExSZwizuDbg4TC1i6BFDo1vgjXq
wV25c1f9rFeR07vV4jRRUfAKBJGu02/mPspgcKaOjuSZ/M5M57YFVuBpckN2oHN9PUg/Ei+Ynbhc
X36pDw4I5tDoLDMYKs5YvLkWGEFdZqyXZeSAemQ/pc/hiMGc2MnE11JFBzY+o/eAPpH4YsIwIiT4
RYP1/YRiHfARmCv8PAe/vGeg2nC6jbrYAAm4UnhE6RVFsk+eUvgjWojcDe+waPK0uXCHeejI9C90
zzK9GXVz9uPqCLJb7mM2XmgNcxTm1tVrxiiMZ4jCk/Cp5O35OLk2EvuSWT7uPZe8UkgI786CwcKZ
vUn6VN3vL2VfwW8dfF6DDGSiJfzaJL5vMFAxuAPbn4tS6qrDuHM1+l8TdK0nU9lf+HrJiJiCBeQI
fzSEtdJAqrgzWJF1uy6FcdnJirqmiMW8eFLFYM94yFqH8ZlQ9fwnulUx0GnvyCJTVf08ggeI11Lj
rf9vF19f5WgzbKUGu/kuxQH14QInHg6kMrg6v9tG2jOPPOhrLzPohMWnKPj8JzANp0WKIrtDZG+O
NgHskIzfmyGqDb2kSDbEgqDqRVjlA6kofLnSECHKbV1Btevju5zm4QlTmQSnjexC1NF8r1BZXpN4
7KuOllnBzzPvtXXVhCp5zwyWEmmIHoO+X1k4Y5PEiXVjw9M42cKeGqOwGDaW3S6tnfAV7J9JOiOJ
MLamdppN/Mlh33eMlHveKonjvwvn9jWuqh6dZp0FdvPWWBhiSI8hOrbfSS8ig2SXpNBAuTu3/fcg
+sTBnlQmtdg6iYJyDG5Q7piSHeFI5mH8q1fXrGRZ+JC8oFdSfq3Ni08IrAgN1lg2HfA2S6MgGahS
yS1JGJWwPxuDJ5ksLrf7+mzo8Otzybptera9skqS89jdxAlwynX2Gk/8nuOUXB3Iqgk2tZgw+GBh
y8ONMe2A59vx1hKQIMJYgybYLprkbAFscijbWckAxrqYaaELGNAcPmftbjdwXVqAFTuqyBIwzH/G
fQuV/wLNmdk7rEGeduhm9Ns4G8mvtwNE3YSwNS+7EdwbMtPPS9pergtm0uTBFhSc0Zb5ycPIbNYZ
t9odxMPej5HrqzerIAjVzMUDpm5xFM+pL6BqYJf2qFcNV9GkYOB4JAv8qAvqa4/BGotizRhRUk16
wt5QZ3gRj60zcD0Fiuo3/QBPnjPiu9LCvXUBFWJQHRfpzC7HWaval5yBOGxEfevUrjCEG3npN7aA
RIJjtgrKQFEyP4f6ABJzMp3QPnr5s5Qkr5Mul6jULxjWRF5Q7sHvG0hroN7QczcK81pdmYjHJMih
jOGUFtwWsRYGjlbfu/Eh9XATrHTFtSQ0VCcBAgOXyaqrXJJa7IJXigIL+bPNTDfNlPnRinIavPXk
NHN8zuWS0kxOZejxdd88HKfxMK4gGDKA9ZYEI9X/EtU22y5DXzWaBrqbAOrM7OlfE10+6SbC42/D
jxsyC3HIKxy6mde1xtJtt/ftL83wtw3u5rkBUFV0bmm9HX8mVJ0z5CB3EgmuxwpE9/OChc04h6rI
IDjPKhtgozDw+XYkkOcu4mNDTXZT7xUrlOLC8ZYDI7Mg7vWYM58eG6CLZLLUCQmL9xZM+GpNv3sv
nWNS7wPcxXdCvhN8kwECgquyKzydhOlPR51xJSXf9Pi1m/jJaZPKzkkfhxi4UQSJQd5wmlfSwbt7
4dKHhfDkWsr6aefwJYCDbaMvdk7fgzwhuECZvkOWJLLtyvE1MtX1FIYjvJ7nc+p0tfi9OpBZnvB3
LXdhE8V/lMJPJFg1bmEqLjy7UqXrHrZCluN5nBgQmU9dk9S6R7waX5+0sFgr16wsCPrKBzBRM1Ne
4IRSNXIkaWLkW8+48yTYcZq6FTbmgK61OnIAMrmoHntEGxwcOo16Q8i1C/PtaGQMwogyHf0jrDcl
AYgDmi49ODZxKy0BNfeAaen/l5pqSn4rACr5IAqkBDI6q1JMrf8/7igUrjJ1J2dcGts+QHaashNp
pQrwlHqCgGSBUDhPMOd98aVD/EIaqNzkwdpytvqhrK9KPKSbV2qLjbx65h1A72qLJaPV2LV87DhZ
jIg0FbG385Roaql/S4UGvpl3BkEqO1ezs5eMb1pNJ0kGCJjxHLm3sk0uc91PhlfPlrydo3uCByyp
Vc2mEWMp85BYuvPcg69zidLm5EKyQTl+tQZmZy584asYxrx2EZNqziuFtkk1iPpkz7YR1f1+GVaF
jfqujtUsXc3vtkzkRZIrlb+a6GowCa0a1ufUXC7yyOG7m5tyaMpEvVruR57qeMeWwnT29aTqVR1P
EV7vwzPBqVvmk7HnzlA53epsNCSGC37kMVnd3LJR6f0i+mkxDJMmVUisux9iwmT5ArLyE26uh7tj
i7wBi2YX798DIKM591xNK1mfOI3XI/NUJaFDzmOLBX3ghN8cP9QmKbujwONXQCfjxLKC/rLIky0w
S5xEuwl29GjqPI34cFn4Ueto8NYXx/UJuebjDPJVFOgcaXMXMHMFUpq9+iCiz8OBteJ0yZF405oZ
VryMBGBKrJ+T5lHX6nl6TK9UQ2M1WYQ0H+mrZzmEwZ/Hz6JCuC37cRtT3ig2tOnU0PKAmKbhtbRh
33WJ5/cvv9ymDDlA3zrr9RMwI0Y3sPmOrRsNB93QQ2FB5RMTUg6J7XfIyM1azmu3psbL9kQsNOsR
8JyJP+n26LxoB/+M3rJj2j/qTe0M14/PPug71nMd6jE9C4c7ZsFYZjKfI+BE2iZ5Fz0MdpzXlOoX
+l8/xG6WtLdy+hx3eyMBgZu6bLidoUFhrILHo+hZ0oxbXlIKOFGwqeBVllqkGbFvVu25wuNXSvuM
+mm858roRNCOC9K9CkKZuuGyz9DRi+dFVtJ0gHhCo80r+P8/Dmp6neDqQ4QnPHnjnOHMlW4kUagn
Lw90/k5YSXJCf4ViZktVIv2LpE7wOx6aCi1bIuCnABv0JDtVNwl3qltf/mMjGws8WvubjJOTbVmX
CV6PD7j1+9RQlq/A6lAaZoHB1FA81Xnrk6YlEr3P4fMJoNes8CrnQxfR6tk2UAYy4btg8NEUpAX+
dXHNLdkIXJNYsVyuTA2xOsfeih0IkR37l4Ek8gQEzcK8tq4BVV6pTvk6Qttp9sKbdLFX1d7M73q6
8onJkgassqJ/3S3ZPFwH8fcBu5ddRF4cmXHYTj2l7SdYSwYpPEgvZO/zztM0hZv3/3yZ/+3PLU5i
tMXyLl0w4WpnYH7gfX8+hY3yT5FUheJBRT9b8LKvdq0SqzY2/gcZiYRaYlhuBZjazyY+vB/Vw6av
dCTgAGFyeuICuAGsnYmBI5BdqEzgrsifCapzXLm9++/gNpg4dRXUD2bkgje1er8Ghprnc1f1VJp6
vv5WDCmUCFemw5i7RxTfkAaQc9IiVSXo4n6Sa8aWiXA86RRn1Ds6xzPYK3fiaopRnjk+M8ms1zVj
N9WXgir/IKEDzadr8yPzT3aBo+7oeUOb8h6htEM6PkCUaB8dfVHeh5Wk7ODAcvtk2EyCG3HxVb6S
Pd89q7u2CCDl1v+S4oOebPVU+MHbYcDYHLU13x1DLk1l0Rxo56AZu/R4UjIrX4BLWpq4fEuWQ+yj
WjVc88dT8ykQo/Cw0gZ+uDpmwUVoVTlDele+e/+7lRofWMriI/FJpp/NgLK2THrQhV75FgW/Bmvu
U5IhqnK9SSP4c5veuedqcAEP1DUtoBfRkkJIwLWOHOZDlAYoPtf71bNl1pDQWIK1nvS4AzQDgpmN
1glO5QhNiYqKVjx36yiXgwpxswvf3FXV5/BeYcs9LRYRZq3O66Frko3yac+Zula9oAqu5DziQ3q2
GPt3xIkTOFWeJnwO/W/WnqR6ycc/2EKa5TVGyh3vbFCh8xEDl/2F1h4e51Hs4tl3Wh6bilcOoe1s
GiLdvTJeBN9Q+WpK/Kq0ExVhDBWfJcqLemvawGy1V9+Gdrj9zEChT+hv9zsYJqkb3Tda9FhM6NF3
Xduf6q6hBIRBFWp1CC15GWIOTJ83FRY0W8gcxVrfDTHa6RdsKJn/JSk+gZMSPqBUuzYL5psEJGXM
y8cqh3nJX2pxXlCA1KaAFixC9Fgp8RC8lWZ1j/LsRN+9TzwIo3ENH2lDcPjho4l2qDJJAjqYgZhQ
Oh6NSgLf9lVL8SVEjpfuDMZ2RnxbvEn/aXRYVHhW6YTG6kWq6AiMdIEPg7VbYnEZY6uhD/fUnjJ8
RAhddz032rq3nIvboNoeOEnBDKnrNsnDDjx1ZqEAHxkKdwQrHLe4YyB+OofXLv/EfSdDKowF6WKk
TKesTlUDp9YxYqeUdN5HWSWP/HtfSFG0ZHJ6t+xmu6pmtZSNjQKRpCvLWjzHBsaTQj0uPM1yXUuB
vJBUkHQK/TOamkSoqLpk8lG+bA16qmfLvfRKGCEtMWvT/fGKPx+6MPyNVO7O1M6T2h5CxNEomc/1
BTAYHnJAD5Dm5LmTaOlWk7gHNuYH3KBSKOxNVoL4V98geRZcjdMVcniXKjapcIamg4LkwR+6CBp6
Pps8dVKWtwRYzilTqV6eUgQyvxuCplEIwUEF2FbLO0+g6Am42LDPuuAb0Z3mIwK8G+DxE3/UOzst
mskM3OO2wQTAj+CjXQ8QfodG1VA5Qt31dEDkCV+z000hNLpLkma9QsNKA+Lh4U0J40ZWobc5DDVS
we8Jj7DReFp4yeIiRzW8jE3cpzFtdWN0SDXVMBrYNRhNAnbrQznut93hXvY+AiqjsIgRLIxrkIBj
rhh7igEKzSYp4lnAkmznYXGI5VCzvFaJiRWedXNJsc34qaH4O0lwE3CXZ9wL3GKpY7D/k9lokTUr
71U47WOiGLgsDKwG2oHvMxzaXj5FYc8Bvts3gnWUH+kdoHwXuqb7pJDxXYWkGzJOly7dvfOga+Eh
5YkveVxU++OwrVXZg7IVur7D8bSizEvUHOHcByPgWUMP2HLP6isoi9q+5eD1spDwI907TT0bp1H9
/DmkG3tvsjWu5lbUMBuoXKCGmeMsvo4v/Ouer9BhFkWCwSUqW6d+zd+gwhGtd3lSjb7ye5oo6WNo
IBZOihb79BFRZ05roWAGocIGBBE/SkAbRnYSLEELSNtCq/2WXZjy7Jlv5rfeCetXbhYVySADzWYF
TtRA8wAeFR9VRgM9yKWBSpy32SncjS59A5misAok3O7dHFtNv5YWk7PZr0SYa4AjtBb1geiHDfou
6G/dI+FuQsrdkoxFDsLrs+v9UgsrKfiNiC1/92BESFpWxqpJeK9nLoxGnX4gs83vgT9B/Lzrq8Tx
V9/I2wD/pUXFLcdtZ+qa271mvOHDAqeotWwahxzxt7Ag4V9eId5upiX0qateOC0pz6hPp8o1NDvC
iPz8MLvZ7U4SisChx6m1+0nqWPXnX3rbcMlbXtjgExkrgaFyWyslHjf25r5T8P1sPfWJ3dbjcYDh
BfPieBVnK1F5VVBq4pkYLkDYgvB3EVrThVmvcF/5h0ENdU6twoqKtumy7UqBQ55Nm8+h2u0BaC/v
KUSL4XdObIVvDTwycunSv0GnVGkcc1/EaojD6UEcCX9Y5YG+8pZvapTHLN1qw+8aad7CjBDDN3Vk
yCxCIBecWEgC4ovS2EJRE4d+v1nXUpVF35fOwLowmhnlixjZ0YwwXt5xWoy43GPgSpQTpxn3Sxrn
lDQ6nl3px8/8XVAy++YtlgUytNM4gDvverK32HGyCOytVvldh0j5f9gnrIL8fhCZSLISZ6ij+ZgB
sF+wPfWN7eHu3dg4nBsNikVUxSIqfHFODgrXCBeaXZZ/jx43+UEFZlxBs/Z6NVwndi/JTcst9A0s
31lUrpzo8X8jbhwYZPakMBX440FdNkbGN7eIlFoeMl1qvCSNLKaWy0//PpWZS6ofCvjB2ZsvzblW
1au9AlrzGAOyy6eVD9pqh+pP92+xP5nk0cYpMpPSuBIrjEQMzHOqMH4bPoMQUdc5HyhLJXuW4uw1
bzcSQNjkaeW0t5kqaCR2syFoFv/NDS5/vaBSaS+0IhxYRGOxQFDPSWPnfPdIF67XRrdgmnC1vKMQ
iT7id9etPb+lgAPu9HwtR3yB90ahXIw8S9XdNkZbjFwapD1atUfxSLhDNpA+9ZAb9ereyxboB6jw
XNWGdFWh9zPmGj4d8KSJyWJIQvaFgSlAR9It+NoH8YjAjXdQvI1u6f8CLwF35ZVKNQz6xNhpWk8A
g9pK89HVhAXmv8qj4YcKzqd2wp8mDjCQPZfLDU/KUnXnk1jjTH66RLLaN155mjx4SMr97kD/HkLj
BZNosM/OFYpMrVkhCTUiPJEda7cpRSVQ6H7ja2nh3raROHIEsBtpoQi0Uq5lgh64RMNwK0Wz3d9i
ST/sZoMfZBh/98Dm942IWXOAqUZF8IZCt3EvTbE0niCyRahTp8EKMKMRJlDDypQQITNR+F8kQtuA
DKqzQjRvuriRxKZFXubcDHiDvt0Rd6WO1ZTgbLk8iGJcHV+qmoXkr2oC97IwmS1HnHYFc24vbusb
Z1uyiyFNlBsarh2W5AntTCHdpRK/a44HPT2VilUdmscsvCSOis76Xznly+Bh14MEXTr1vT9oJmzl
7WR3E8zYya+HEzoBkfgNbVwUGwI7Z4zO2t01LFjg2ErDbtigLMrVGzrmB1v0q1AfZKD5zj6ZLRgN
2/Xv5ssqvSzBZXqkbNzgFF5aR6c/3ux0yaceACdgZSe390EWvabaPk8U12DquGKbP+cM/ZDhwOlt
z6ccVqOblwxG/0EcjaztcAyKe4Turl/K+9uHwDdirhs7U/oKeO6mV0Nt7F3cZHZAFemgtdWfJOW9
3s3YgwvXRzGfdvXDqM6CxumnFV/6NCDqd7fEH3i54+HkK4ZPFmBjjW17Ptc8U38G4M0ZSSYZi5Gv
8uxP4XBy2qIFAgzmOEvKgcqfVxz0jp9APUJ6WTJFTNOvP3ZeHUcdHj1y+J8/uYKG0N4T8pW+Wem7
Ax+nRjtJ2Sueiyppcy+DQFgLFlE/sJo8EK31hKb5JPLHOBQO1eOytJvQqjCBrvXR2V/YjVp+Z9ID
/5RJN7nLsgzJuOZyg6ZNglf2bIQ7XasSMhQtGvOZXVIC/2tzGt3yLvMmkYeKd8Z9LlCQhRhGeOj6
szZVJ4tOQEs9vl3QU7yMIB9TcdLi6ctdMTqfHkyDK/85TKmjcgAxKE2FLDeb9+tTkxnxe52yH9CR
a9Z039d3VtD4Z52eEeIchA31ZSVL/dXQzUmE8cqdFdE50Yu+6e5DfsiBbN74WVExDiS3gu2ObEQc
4GDEo4zoRzlRSgpwkBSDKR+sAt2dakoaaESNyBOGj2MA1C1V8yl94gS5R6/1fJqYDP+0brfY43YF
RO2QWY97PdX5oEGscleBcxc4Cy5KdfQ3W6k/tVdDLBX3/zb7SOZnO5hTP0qVFNddNbxwSMj4ENHr
kud78QrQDSkHu9LFneOjWdlM3VzGYIXg8h0PxK7Zs+kRlfmW5PCN21RU2LqJK/0G8BYJDFK9W37U
mdVTMyAYfFiIqkVpeG2jhW3q2GNiqCZHgEHkkJTtyQrcmG2LCrqiDA6q7ZpCXpUPN4Dy3yplRzz5
Mi/87pWWSFG8Rr+5F73kZPKoysexVOszqBmnB9KyTmqmGZBI3SnsZtetPxkS4Aews7MdVr9mcOsl
kNhABWjKKp3IgqpZvZHWSbQE+B07/2dDoRFpw5cB9dzShoOKW1Gx9WzfnHCcp+6V9QpGEm+9TWRF
tRi97MH7aBK1c1uCwdJELlmpZLnJlwjksCNP4QTzRo0ohZ+lGVNpAohMnBQLtmrBjvPxTP2/2Ecz
UwxDMbX9uX7wUBQQbmZ7f26EMRZbNwro/eWwRoS7jlUeXVFe2RUCe5F+IH3B2yY5ngzqnfBHwzfv
TP9KG7Ap5eEcDNq+xDmSbKCbbyYgece+bLJEopadgO1mn3o1x7zoQ4KO6Zy5Zgxv1RSyj/DcjOb2
vCJ6TQjSGC5IeIYF/XwobRvUaBVF8AKr9Zh3pSiGqotCy9L4qhmHYvG3sKiIX5XtYB3Ld6hwiX98
LLYuUAKvFtgrV7ECZmQmaob0R9LpPBf9pMgHBn07XEGrps5Mex2u9Mm8lGRPuE3TLduXHhXype2P
Imp1pYicvBs0cnxImx4Tvhj7HemeYw8159KuGQnAZ55wURzp01bCBznm0nQqTXXaL6oz7ixLqQgh
Reb9W4FwjOuqIuZajBF+OXzbbMXMK5Oi52vgbFRbep1MjKO3w9Rx1V1v8Ohhks3a+7gUqaeoKHqE
Pb7krGkL/PAgpCbgJhbtoLXPlysGiZftit1nkoE1c2o++dAcl7hKbvEIX+rYLqBAR1wBof/0Ajw7
MUie+CARXlTtsXHiSTNZ/r2eTVQY/eB5aJUYeem+VGAgeHYWmVmTjB88uL0M429Ae4ELwDXxSQJI
zwp+S/I1fAq89VWcAqn1EztmvVgcScaJaVM6cjcAll2COie/mveyhSEXytorIX84jm68jCT4MprK
04toaubA9ORHUcXZchJo3RlzFWh5goqD9jbRC0GMtMOv61W3qkPK2PSn6l0VGSu4AcISkQ52N1xU
4W4RMNgfUulVfmqoxHK1d7mVtaOFyRmzH0VNYZguAxQyDDWGmse22iDNHDoLhBOfrJL26pN/Bb50
g5A31P+p/QI7xswg6dFZD1ehB/51NnVefS19hus0wnLoGtuMPanxdlTYnt6WXxJpdlVQ9HV+TFzf
QIm1Hfk9zGp5b1yOnCPcMWjKDA2ZpN94Y48Qdf9dIpJ+nDiXj1fll3llcn+UiZ3ivS2yKHVqwzpF
x/uakqWHwcPjRkUUtwUfjcrvjF0sk+fzwoib2kSpAZLkWMjg4iCsM4WW7j2uU0OSdfxS6he3xI9K
2R5gXFYlATTc++vUXcoDBc8OarMIbymdxTQExPXq1DlT1q3yLkovpabRrn8h6cM4Vo14z36G4RBt
ezLo15hg8t5bnqHJCOTopRXSir1EodSprPr2ochSvhXFMq5AwZg76i4r/qagTHvD29x+rXC8KsR3
PJlfXba1swTGaensCo09yulkI9IeqRCu3Qe5vMsDdZ9J6/BamGdlOoUWAWH2QhcNLfI/RAaP2RmZ
pqkqkMyg7cS5tZAC4BdU5+NCGsUU+bpfvdDH3HEG/xi9aX9jd8ONJputnLXETsE5eQAvGn1frCQY
w3fXh3Q66C51bUev+f5BVQN9TY37No60ag114RA/apfXTwE14vYaCtcZDElYCQsnhhXKhc/vIofH
+IE5kFGc6HR2NVe285nWcZN78Z2Y5vz957m7ms1wRMI5inNeOtZnneI9Q6A/mzsR2pDKTntJfshC
3wQmJG3SuoGkuAD4INTFO8nfY698sAI4EPLelja6Owgkx4PbtgB9vUQ6KqzhGQXjHH/RI2/adDCo
I7Sis9e3ZTtpjE4vOeLas40PFpC5p/hesfYsv8bq06RBuJBjHL9KL90tkrFYgFDQYW/Ns+j2YVAc
DuTNJ1u7O0IuKSKhkHV2w2U6dxtZnk8r/Ml5MayFt38T4Uf5P6B2f39JEC7B8YwnAcKITq/RaFBf
7ANpXAuMow+hn/UFXfDI5JaZg845drspNNSTo5fUG1c7lAV4LDKoE7R98pkCQXQab+YhqdRp9loy
bSWODy+QKRc2fUWieOcVkeKpA471dWacQvGrUKkOeLXVmAGAjBQJz122o4uy8foCXT5zQ1eXtyRC
qo5KAaEhdAb/91oNtBmFmDbX3LiLaEVO0t2lTIZH6h/VWNEshTri83bmaEkr/8JEwvg4N2tYJpE3
HUIWW9zTn50OuRYyGM8860Iul8Gd0oXL3I9KfNSvKUd/9HI5ibcJ2gxH+yGTtNml3LDba+TYV/Rh
Mn6v1IwPoa7z1PgAzFDHvMgXmjwBR9VT3d8mhfvd4HkDidr4D+f4bVOJhjFFazooM101/RLUZqHL
pU+R0lBm/EDekMj51OnA0G6P5fGhugTdpRmr9hTfYEtd7FmXDQGvjcWp1/ahyb9hwAF6REVtFd0P
oPyj0CDiIJZw3wIE56ZnEJhF9pVGp3kQWJtU5uuqdd4DmIeH2zYkI8Ycj8CQDrIeHJJCtMQW1JO+
oqehQT2Br82A6x1ZaC333P/LU9I4bXScr8YOhar75p4pYsztUVnWIuCB146MRjaz0Deb8YRTnfDn
4RtR4S0bvQMFNHBIeO0I11zzHIG5f3Zoz8k2uCIWjQpgi8HMEFeuK2yWL3lpxWS5It7SuuiBzHWo
LchwoB1GwNLzFNULsl7sp4YkV28a3jDtOfFblQlRk+sv0KpaLsd3+/bI9HrGrskXk1xivwXDO7n2
TgfrXqgr+isAGbANBC0yTNcH1rtUt/3NyULJDFYT04LZRpLEigKlJrkNHGOLBqVpKn3e5junYMT4
wOqzRI4sjiRo4ilho6x/Tjv6Sw7HsXSnwR92pukwT1YYwLyTLwpZC6ZbaDfVaKSB0+Mk6RhNMQzd
pZlAnH7/V93c5FTkU3iGhTAlIROlJWYWxrB5m+S2Gl9flqkYHBY8zX+ygW1XHIqtqcTmwcwbRUam
dF3DueW917w0ZE2yza37HnqzusLVX8FQG0IX3fQigzYeIM9kpOeZZQ5ZXSO0fqVmOM3N+hXXw7c0
LaaP6kN0A9bxT1+PeOnc7yNTAnDDbs2AnUP5eqplad1JxlDRJsgKKEzP+R2sZg7FATi6hkLDblL7
DKbQ4W/L7JvbQmk1E+ka/jkeC14wDW76TyJEfrqQlrBwHA5DHc8MiNwrH/MANAFruz7hnJ+IbdoC
Re9A+55uneOKfwlf9gpXM+RDxoJCUdAS7ME5VbJ+LsftOD5H9GsjFylNzb4DNXB4wN806cx7EiH8
JbHnSzuv8cfiMu4LSMLdJi0zW8aBjLmXu38wrmAdvIdxIhATuN/YxmI4dhD1QxARV0YTN35yaDko
uRyxECah1i3uxDXespPOmjeTyEqvD7ibI0f9kN9VbLycfu4sOat93HjovBFsDUO5G0qyN6Pq4vAG
0m4YDQXeun/HOAdM+zFPbxZ1Q/pvbQA3ubj4L8u9qGyLkhyxaZJbG32jOwZx2FKMF9Oy308rJhE/
n4Ta6njf/q+3yJq+kLNtNt6l/k9OoywL50tBLRNkUBxMupgdS0O2tvs5yCNPBMSdxhtNEhSLm3if
9IuKw7z+cs545NoPeWm8sXMHVPFdcY7oGXZeYISAtiaPsyePedlog8GPUZlLcuQlYVA4I+G7oj/O
AKuyCT7qIFAadkb6q0XHFB2/2vIkVQweu8zTrvfk0KeUzsjDXUWv9IogXCOPP66umN0mfwaWtdyo
vHrTZMKwUwBqWul4zeWcqUQMhCA93IhfCEFNjvdu4Zr4B1cCtsH1mSFX9hnLw+YyUtyxPF0ZXYJi
CwwBZpp1QhnQYyzjf6CIu5PTUNdebtFpx2HhGzIevNOUBv1h5FDV5ONy5oCJvKKpVfCw6AJnwPal
/RrcEldDH1noyf3dXosIr3NqSHaPYyAz1niCWgL4REgsf2/vlRiUj2XTNqVxBebNcuamHq5wXyFP
3l8hbE264uNuLFZFxofoG2V0usjyc6EM49tjsx/XhND4jV5N4gHe/AFxKKDK/PQvzC8HnpMzJvnK
q+vbjMlUPj7nMCsbLJ9N6WHL6KruO6YSUvpHxWHvQrOJa4FpGzfLfKQbP+sU9MnanB0EteBVfC7e
RMas9Ybm1TI7j3pAoYP0JW4gBwP0tuvvTRGQO9JKNz/pB6E9seN8noHdYFiPdnJ1VWMVPguPA2n2
y5tolxmP4y5RTEMVgLGD5U2C+FxZkeLY9Srt9HUrffBEQlh1f6TgzKuKETPVBTfjpdd8pMCY/YvV
LUF7rhqziKEUdAnpbN2b3Mwo606HASSpcKXWiTeo7ZqmousOrxnfpa5s+ExmQjtOkS+11Of84Bnr
C7+RoLSIKuwxGdgIr5s3dEOGb3lYKj8dhcozt7Vi8i5X9lCIBfD7Rj4SnvI0yw4yCf+PPFlcRHJs
EqtQ2BsU2oaJHnsBhsKTzI1K0/HgjbSVSMaiSig718f01uHWBemFrJBLgQiXiCAekk7CjZggD6/h
3U52vZapDV7uay7YswpLO7PnZHwh7qLJcXVWenWselizUB049jCLAV5x3Qgv8ZJJXWJkBhbVjEPv
4v/cPrrTc7IZEupDxzG2ItXfTKP+8JRaAnHSl5eiaGxF+IXlTG0DmATIBGdjhFzl8LBeyxy42K5v
n/V/U6Hqi8Yhru5M50HGTwa1UjSoJOM8Xux/Ll4R9GYG4TBzw1IqUlt8qq0QTKzdJXwQD9rprOZA
0dy51mU82k0r6g3ut+EbMt58cYyYYyndZi4RaWG5rBy1Ue3ZMMEOjt96Yj9Ws/RKpTk79LDK2CIk
A5s1eKx6189VJl7VCM3QKGb0YmsLYD8adISUpU+GMIKUNRttnbWqGGymmh/r+gRTYKSpjTFURaSu
moY0JM3lMT+uI5oe1aA40vl0g24/MX7hsjUyZGC2GKso1a/2Zve71aaUk7dxvD3fNSxjKkndRjj3
yvWgtmA/HypqCCAC3yfFSlwRG/LNxZ3CTLK7MX32PURqGGMT7p6VRLv6jNnaD6OD8nOTELoLhsIl
bUVjjCmIJbCrbZY/DP9iWkkVQTDT/MRRA7hWCJkCFXsQ9Mwv1f/1PCBLx7nfpILC6etAADVBqhmI
Eg35px2Iukkm+XehEagsG8r1ZBJLQFW9U0aQtmhQP7m7A3jNDi6OCxQKoMr6Wd/rym6oWqrvzLcu
QpqF/PDxucwjb/GEDYVwEuz+EAgMF9vHGJUXsKFj6fD+Xrk9QwbbxUWt9nKjw5EQMYcIXXROMowD
ximJOiO3ai0biY/VMEA8jBeTqlPcg0dC7ciNbdoWnv34h2rsKT8Koj7cgIKGtfssGX0BAz489eDz
QgI6Dj1eoPVoWYb+/h13caULQtQpgZtL/xSPnlZDTznT6w0gWB9l14h43RaQ8rEnsfuajYUbfUY0
Ko8d0qtAZIKYDQUpziBHpOS3juYO7HkmPjxVqFUZv5ZGRCXK6iT/ezVu3E6o2QzeK1FZ7P9M7MKR
gS3//iWpWNHPDputg+vBpYV7z+iVaYVjl3LU5meR0SSQecWKgmXXM/ydy/FgESGTrZ0ksXTz+KJ8
P2zAe+4BBzSzoCRjr8m9S8SJ4Gv2VbKS0XXW64PXrfBs47V24FVGB66ZEEPfd8raORGXPSpa6ifB
d9Igtz+Xn2t+0SQHr8bccOi9n1ZhHOKeERzPb8DKK+jSmy53MJ65xfCzyeXIeUlRiwjt189vLVOt
HM2ZJ5za2kmqeZD8a5Ic5jQRdMt8SLi/nl2hjuM1+6vIS9V7c/XjEaMXT4muL6qQCe6xOILLzOvE
nQRmjsVjLdfmbvEi9xZ6m+DLx0WefoXGNIuB9qkIfkUkPKLf1KSkXvgr2s/V5HFCvG/8lbJZWtAK
9VMGvEkbiyQUcsl2z38KZGwZq4GQfyxvbI8qDLF/pdthwQ3oN+UAmjmGLkHxAGQ7NlE+q4XchL5j
99PLf0l4NFrwQxwyaAvvWLAWgOKm/v6tJ7aosBrUh5UvX7W0K3/KWtISIOvFNpCxVsQCjVJL4x6O
xGHzgnFKMXp17/H1gxtTXfY2YjS8YMxoOtD6p2VkIVWpfwklrD9MARsayQdYyVYUR6+RAjXZ0XYa
EIyofUSHo6hMf88mcqKzV02EVpcFWHpt3ykCj6kyzNCvpa8aqhm0YZMns9xFzQZ2Iz4Ob/8uiWNd
WR2YfBwEQznEAOB7h6mgaQrjQD1oG74PcWncEIODLBqh5dvxHj3k/VyqQIfI+HfbXCu9Y8sv996T
kZC0qUM4FZYyVpaKVvri+eAh1rLmJidA5hFiiMd7fGE58tFqkA2K10g1fltxuewgwS7M0Zm/rDxY
gElziD4iskA4gbzZtrGFP8hkBKdQHAQZlK9nd7rY++QANqor70Wr5KOu7VtoP/fXfEg4f/0gQPkJ
aOPdx6ok3YFQQr1FledToCmXd/llWoJhgal2+IQVanVCjESiA41VxPf4S4WpMULahk+T/8lAd53o
Smd9Ov1dIGoi+zgxxb6TMT+wEXDm9ZIaE/Q1L7EFTYIUo9i7fXJktslwA9kkOoJLq3IvfXrJ7s2a
xrvRT/863AgJeG8aNjysFZCDGrC+WyVxGSXlojXXTHwh4xPvaCglTEla7Ttd+5wAShrD7e9VXu88
icUiHKMSO6XZYobKigE7fCeLmoy16DaFrhFIjwAVUsQqHPW7N/bTXore+ji92xdIam3PzqB5nIdf
VwPLb0vjZ7qvnER3e9z1QDexMI2RiBgvVRXjDNWxabqI+vxapMjqbb6ohSNwIU2Idcs7lvyXDg0W
dCCWhyMejox44SzSMs42Hf76fX21cLVrIdd5j9rZ5Cbuj/ABsZXFV0nx9mf4ORDmQUMuZPiqlnY7
g+kkNIuIg8Nm1yjJ97AKtsWPpkUxitx8h+56jO7mSpi8+nHtjOCvAjHX+ltQdsUMv+LhF5NJnlHL
0JDeN5sDs/t9jc4mdUu1w9J2vsZfJ1FmTrRgXTxcbqynzi2/pmACc24zfp10YMBsE/UE8ER3hjm0
9TUpSfGNH6vjyBUmzQwGjcECLf0/abFD15t5gD59HbFUI3wocPwPooNy6YVWEsk0DkZR6mBtYUl3
a+D4tMWD3Vzfs3aGa6cl8MMXgBo3L84wEqduFh8i9oj1URPgl/bzkIzf9KKmeOFhsWbx3wjvWQPd
DLVV3K/j6WX3Ls9vQfSDTxLIjBCGbwdnBSFMXkc811dZ51LFuCWoo6/ZN3uP+TVMh+pk4PhanM7W
71fDeqRxHmsfovnkzc35atcwe+XU4rzObNUxWzZ5FLG7WRav2CVgK4fvtUBrqFIo4LjwCmNYMudP
LvM0i6X4LJdQgwzo7seS0JYTFHtjmMmoom2EbstD7ZHg96PEf6FX/UkCu6dhxtom2Dk1EI0upPOT
U3VBtRkg6BeBv2/nTGFyZRVtwaw5E1tt8GnvzF1ITW9nrchG13cpJSPScxEHq6vaI6fw5s1biwqs
NvtqK7bzXwKT7mmKgIZQ1sUbWDN82UFpAHYvsA+LBZ/yYSDmZeIHLw8y0eQtAxC+/kH7/MGpOAhI
GMlahSSaOcAOb/XRlw7aVPT/UkaVMo1HaRMI1tIKCKb58FQ8K5Xsnf0MZX8/Yxjz37g1564i0Kze
iaQxShKDSfl9Ly7dnhdTco8Z7RPJTsoDPpzeqQVX3BlGh6Jocw+e4AIEaXKPoDlWgbOwg5RiqA1u
GN+Ej5VGj8qLqIuJaEBNaqEw8Us1y5n4PnHglMM1r827HgyrHDn1M/Dp3QjNBgH0WHm4Awerq6Pe
XTBrTwyVIQQEaeHBCbX/3BIluNpE84gEU/JLDxXZMympQrgv8Y5QnzgiCx6og7E81aFuiLFepuGj
dgPHFi+i1DJOA7RPQvBUaS2k1vDrLDBvmw7XbJxgFf1gMCPCPvmviugPkTSrzepaLuMhajIdbmi9
TXiiNuKsyLH+Rn3+feSXk04zLJIYfmxR0ksTYY0KjczYqWNJb7CGSDaDXMv6s180z7x/1KUTtkdz
2Nw8Q5b3f3Tf1f9ewUdhTX5vXnsQcfRTsWTZ5UPpv3xpJJsUzQbZSvRCcIE+BNGo5gwG8lO4KU0i
8iCqrKwzDKdMVtq1EnpeJAYT4QYs5L2tDZZblnE8vwArQvFuj0XrnR+MBCKepljcSqkW2mZbkyQq
vTNfzupQS5IshSz/DmXjSzk5Pdk9wISjPg0bAgZCUJmIn5ePyuLUadKOJiVtwSjJf/Zl3b6G56Pk
ELohMYw72zjFVsVPGxkf9WFbnptMWjO7hfSTPE5zwji/9bV1rqBQB8OZ78ba+6OYCrY8nutdV8ga
ZGZWGa8bCigR2uNZWEfWyfZERb/fM9yMf4iKgelOuIEzoTrLrra5il88gyeQBH65mRGLqI7Bf0b1
IVZbPVxoFLKU65fSROJnd6M8A5NqC6On4vQxNJldbYR9Zc54fxVi8oAWPJsnt3DuO+LOAJpRHCC5
J9Ii614pASaQKrVsLDeCAqVa+a4ttXKuvgxGQetlwElnCo1apNuKzj5PVOSU2MwItGzgXwqU6JZm
U2Aa87t+HVjluUUAZgkmZj8ucXEt2lMK+1QR846Wl3HlnQJbk/XaQr+N3CWqYHEsRkCwMaXS0spG
JQa9nzIRwcEeQsOjenrZYQuHP+koUP1O0hiGDMe9slJBo5fEb2NAcz91jvzRyJZlyVQ1vounnY4z
Hh7HgttkbSxnyYxVeSVHNtKyR89kfOQh2oEgR4isB3cyM/rRS7tmqpTAzooQ2iszk1zo0l4P0eAf
I7uL6ZiBvRFGvapgMPDTtE6WFJRPmK+E8xPrv9phx/DGdcYfN+s3n+hLUbMfZ1wSvHBp0TlNEzYp
OyCYnrcyGngN/hxK4g5HpZzz0QQ26bUoPDFzlhsp9+pZG6pqwxndjrDVQSelEul0DZn5sN6bsMlp
SyfdH07ONJd94FxbaFOyrkCALQT8JZI6E4OW1HoNmzYJ8dbsMn4oGLYp1v2rT4Pi+6zouC8TlL0e
zoIC+bXtvagpPJKw9N40G2C3e9u+WNPgmcM4jGV69ALtBd/y/k0dse66XX3n+CWtLvMnkBFSWV36
hfvafHbn3N+LbIK4JvG9AvWLUcmV7D71QcQPKAMHNTBaWJpzcYL0O6YYi0deVAglQn3R7UsN5vo/
kwYBEzT6TgOYxSTvPHKnQWPwcwG8xoq/TImrBKEOCZLxYg9sbNQz+euMOEvgiD//9kMpFKyS2rDP
GDcqAQ3ghmcNBO6iaBQhGZ1fhlLA4syTQH9c2wrHxjTsSI9XgApCMzjRe5qrw6q2fKJcuznmeWVy
Jiawx7nO7l+KoCV1fkOZj9ykzs3bCuPLfaSoXo6bqyzuULkqhsqzn9czA62+O6xZ2LunlDebl5UV
ZR3O6X2hupPGCUpVw3EoVNfTSgZVTYceYgOqU7j+1l6/DLRk9ZxguBQeWFjuKe4M6boqW/urf/jq
ex6rRxt2TnvkHjrOPcQD/LGJvG06t8dMTeYllPIcRj6f3S4p44X2OCyIYr69Q7WcclrjQ9MhsVgU
eLiEPpXtkfQlxGC76qUERPrfzUccCKM5X+gLQIpo9vfLmHYGj0uqOfEkR5CzlpkPEtdFo1M2V2dd
V+hrbWQwOQrfpoeZ2T8xh+qGuJwO8aGf2jV6mVmWK4ZKq+bp7uL9qFFt7tNAEKKiMnGV7LMP1kQs
9LA8yiMRPFMNhN0NAD1f9YuuiF+baVrQZ3njja81oU5f4bj7Z9XrSr9OLkmWQjf1QtXo7F5x/M42
o/mdNWF8D99785wrIe5HCdL2QkBvYZAJC9YrtS3VaS5CCQpMX37ay4MnjSuMdGnJOIxjw6edk3IC
bsWxg41RkjnkA7fLx8+hg+WI0PQ2kEWLaZ87y8O+/ehDsbywvlQESXrb0z/Ai5kFWs7e9q3cr04g
ahnf53omNXCnexgwSmjoC+CoApDqlcje0e7IH7rbKYoJsdB1dTZLwSLI98IZI1RJYfFpz/8TRCeO
ytnvxzcjjQRuu+PfXeqEWQSiNOqa6ipBn14T9sDSUR3N4NMKlPYVs+RMRrGcARVG14BGBGyFo5fV
WeoLRlGbjgXygph/TIwWbblcS0oXLebM+TtJG8d+uvCLMBNji1rxpHHNpqRWMwIXowRsrg9gamRe
zj+Fig0+fzQ6KX+NL6OStLN8v1ejycysiFog7WZEbLTq9gUV8Ozbts7nUolePSZ2evHW6Niew9WY
cg+JxnN4ZW14+D6bHNltJsnAucVqLoR7VqGOwqlG8mV0DWITqDYn5iGZYz9Jrka5Kc9SsQ6YUHhY
DutZkrKpbdHaF8X5W/q/iaHlVXEQF9sixdR1kpy9gI7LRuSFd2kr9PYxQeOaZz//NNOFj7VVLhvE
i2FqiGe4CijwvX+NtqmLR8YKMmUl6a3k0d2QHsJF188SiObiPECMG7mpna88r+Q9hqmNQGI//ZtW
e7hoOvHDhsr1mLictbrjv5BqEjdyg5u9y5X86QRgnrWB+NNvG+R1t+OaVnpi78LalaryjwlmEv7P
3d9wQFkwLhbiz1GIMLQqOm2hIKVreLYmsxUGYkbPqQi3/L5414zHWWIdNf6pPgLbmKtzx4CwKWMY
2nXWsCC+KF/Sq11hJrQEkenRTTpwdjee+QNRDhaIMeRLLboy5xmJoMxRxO1WNtXA9zSQHjziXa45
P6zZ4x51bgNZtpitxaC7yQi39tWHDOI8Uhg7CV4+uxvcX86KlmL5FfddLBc3RLNTzFwWHfw4pARt
clwcDEQ5sQ9apKH9k9M6vx/Xf1AjBT+/AKJBkMiRjVnt9sVl0Qkro28q0xPgGI7CnHn0w3U41jNP
LxS2VQ31JIE97tB7b19oxE8vVTcPEJi+fK67RpBH3R97t0ZJTPoVm95SSIn+BAAUoAYchgrFob1Z
EYeYJJcrRGKJgf+J4SmNwW0Z9zUlRKgWjyJZDnaF0Crl4D8ePtFW9fgD0zReptvtHs/Wh0hrKBW/
1F/9djCgdK6J8vmY37QF1r6fNSaSzlMcnHwV6DYFlIFFT8kYBMb6xmV20aJJIsaHrq4XBJPCoXaO
jSsW1YVeQaLNB5coqqk2iQqn827eszvg+yV5tSCm1JNQnrhwOjbVHDrE9Tsbnsnt2AWGi/nsJW6m
T1eYmxahQX9Dh/J8YKi0Yk+lwaiO6v8l0tJxt3PpWtdwWbrsL38j5RHMQ0eT3QBzG8VKUwZsfrhQ
sUFZ469Dbc4AFZS0SNrFxPMHyRhWq2wQEZ5xeCee3jyVyqJZNz+c5UVDgAQKyQN1hEQkGaaJs0mh
9ctYP6AzHq8nlpmGd/zRaVTMgh7yU3FeqK2/NyjGWF15UKjxchlrf7FpkZHof0beiBiprBawF/vo
HoMPWrQl3ror4OFMknrrvzuz0q1QlrEj8IXViI6q4bgIL2i7YOmolR5zwcTDk4XjTgNQ454Cu8Wz
6INovRF+QF0nwOqiRI27Ij4P6GBqw/BjwFUqL2qpCcTuSQd06Qejt29mbYYAcBdYwzAwVe2kbv4b
fPxN1TTfUeJ1nxZVrRoZUnB1K7xtdLBcuQO1sJSbCg+Ugyf6O8rIYzARBgmRR5S9187NpAX6OocV
/arkJtYRRdjjUOXEmyyU+NOSdkMOdmcYqYxYQCOnp2aPP9v2pfBhC4z/CMefM5ciaCfHE8mNI1hl
txrEH84vz1juwwaTHIvB5eTP7Yi/MINlYM1staj1ysqEZyXXiCmPvk2FrFNmozJus/vIaOWTREk5
L4yXJiUjn6SmeLBqBSTO+QZ/IzWsNaR5OQLv02i7QgYu5av5t263pU53Nv5dJjF80WIKKJYdvLtW
zkIOdr0JJ95k07Fd9rvdYeCgWQWcmm/98Xtnr2Cp86Kn0Fa0m15cFFzBU5xO2+e4f42zgqSwqBcf
rHzOapE5XMerVwkPbWsx5os4JYYzLSFP4xA/ulNCaOvJ4TQJ3Kh+IBoUVmA4Dg/Sbxl4yGkSPp2D
5O1a/Onf8/hh1iCaJ0NWl9Le264qk7UfLfIlhAHzhq11QZ5S2hSlNcTVKO0rd/jBb3hdaYG/aMIj
rQ66+O+h+hlPbKl5JVq6dk4+nZ+HNU6w/oUNroGUY3yX6eqiy+h9TFMjag4JpDb3K9WommkNdwar
kLlV+a4Xr5EVEi5tApyIqKr15ejv/l1ZMWHI7S5ERZfNoh8MCg0QZ9QRZBJJwSBOzSlAvgWB+db3
Zf2iDU1ESYqfBCs3cyhOmYUXZwfSfSmQ2W4rO2WjzlsiGAjw5/mao1o+/61sl+XKMpEF75bcTOpd
IS85dyNXfKiC/Q44yvR6dqoponujvecQu//dxGXwu3+y8HDwnPSl6VkqyWdtYh/1tOheY68ocK+M
2oOdKPsBxf4rKPDcYtULmrJGkwzzWauLJdH8/3kGa5HAE7s9XmIjfQNcHXxyDSkSYh0DKkNfPE8l
gEokoFplfKUetJEHjP7e3Spn/3lqhGECjrSYyArlJigDpBAnb9xDDPIYBeO2boViQFqm7JcqwjFa
OPuTutXzlBkBs/1SlQtA84DrkkkVEhin+zG+PSg/8x4mMcNSizucGQzH6bA08UCSHqDue7VgIeGb
1N7jjt/+Gx1sGtQddWU3fCFIrSxqUHlsuZREOIHJ7BtOxwepmgycqSZqnLb+U3KnmCOA19XRmjcs
YliI9G7awTZhxwJmrWRfYywgEV2k5hcAj7xdQcINrrR1SqnsX15/BbdDBELk+S/pM8eSxKyxdeIE
O19iEVHAgX22zfhRlVhym5oRZOCji6Gm+tdvIf6DHoU0mQRNKZRcOp1GuAOG5wL42A8z1Zzb8MCb
qOJHLjLDXF52PjWK00aZ60cwibA5NfU8tCD7j7d1Yns+nrzjEWprM44m7/jZwZmzTvrqnLSTuQeU
OiiVqCdXyyOD+TIr60Mh7wN5wMjRN28D1BLaXJqtd1tpTrwDCcFd8tso+UxNKGNi0urRP8hDoVXw
vR676BJY616UZ/1cmpSfpDDx95ZfaRwhYwk4+nvX+qKil9A3GwJdr5hz7h9eseQY2qlsk+YfF5+U
CmTdVcJp9lk+d41XSUW7lDcviKpARX0FK9d3Gatge4ZtQqG1CESW3lQVyYlOY1QqZigKjXcLkrb5
+arKG+fw5rgmRRBpxZ2rZyZneIzBc6fAifDPMnNkowFFRcT3cIuD7VNQkKkDrlSRZCrz0TP4H8HA
5S09goCHdWD7Paim2qzGYJ+rkbvCGtHzU+mzs3BQoBE051mqJDPEQ1mOp0jlBBBNSFQ+Vy7BOc34
alpbd8ZtM8hH2k5SdZhFcO3NAJYVvTRbhABzQav7mZKsAVzVAhJvt0/P2s97PwfF7Md3lLckwutG
hWcMWDdl2eckRstk+efvK7Ssn7mKUGAWV6LgCQ9kCzCGJSar6NnWPuzcgfY3nr3CeHMWHDnCIYWp
/F84ORdPPg+t3f8aNSbr6qMsXqryqBt8pyOVaOmHWPlU6ZlqtR77kBbXd70Yzvl/6j6pVZpbOQ3c
2S1OEvDwPZ/5t8ZHgiwRWCdvDNHdDoDm9jhvf3p8pg41+047bleq9SDoa6MUJMwHD1ecVth+aw1I
QkNuCbiobLNdFQHv/iRo2Rq5GyhIn8HTW8iVEBKvJGt70829oMrYQgOM0aWmUnbHWgtcR4u+65nu
1ysXmzqjc7OYBBUabfGgRZjnb3F1CoPP7+eoN1eVqxxwO9MYEY//tU64cPeNstAtS8HMfmoFN1lm
M+GrY0MSktdTIGY5IxVW4WbFW7HOOHqGYYhiaRhNOTHZvROG7beR5O/SVuy3NUmKEtwmWDXvS+Zs
uOBth9yytiQk9/jFjPidn5o9UCNzBz8dzZIXx3wulNKdvbnsKel7C2hKkberw5OuuIVamVaua/l/
bxj2BIZJa/Z80mzWabi++5Mib5WDoPF74Xzail8qzg0XseDzcARqeOkUsht5e7+ceVxq6A0QyIux
tceYvSbOR8r3/Vn7/2GIfx9RyxhiSbDKPBkeCWQ5d/sMMCEEIs/IOo8FdoR6JAIyyVjiUPOerasW
WoGkagpOzWRUll6/ieHmmyoDZ6duqIU9KRkGyeOvP596Wn9GePEt4OdMXkF/UMaAX0Cm44Vd/2FV
CdIk/583Cg8hU1IHGJ7ySlT/5/sCCXXdANeenL1X2MfMQKI+3hv1EHSMmY2ekNULKKM+xA2Nla48
X+fySHJrcyylxq30IrEqY/64xU5khbdVtlsUzsLjsV+90thFnPHdEE4gkmOQZWZojPTXDzs9CH13
u2L31xuziq9Wf8M14Ft/dTe3a4uolFZvOahpQlFv5VG9fJ6Xhn01aRmF2uls9nvwT+8juRtXNUF4
pL0bmXY7xHuuRgk1H+xEtcj5Z8Y9uwKI8XJQtXTzqd1WwEF9fayU+Wc4Ugi2DD1wjY8HTVRN73Jw
5RaHu1tHtQzTBA3KUy40F6SBXJL4YJNsmJ4NuIZX1cxboKIKykX35E2ZFdVQIGYqsWdWijeBX7fr
j440ggyFJyda7Lauej1DOsiF5UWc0pmWOE8ur+gVJ3MS3coBs5IXig6uhHXbn9E6RPZej9+jDQq2
l9/WGK738CHbYGxpgbssC5Vxztn8zTZdCE8pyYHwpieMQZagc9x6H0AwGmDAaJpMcTWFqjCZhgLJ
uyaIVHklQVk2NS5O2A/EZFUhVxgNl9wUDdTTWM0hT0wygrZBgpHu8HkhJyS2t5Ek0buW9NeNo0KT
F0IFxuMWV3AyEYcRNaFg70ORLCCX+PEuoNBW+THdfZcxSLGghzzCqzF49C5UwPNkaimj4dJsDviV
0lYccRrQWUFEvzZMQnY2107cYY0ygHHcI1pmjm5rbxNRwiPH6OnR3seuK7lsBhEjSuN+8PmJGYXR
sHn+R0beAmIvV0ERFHyotaIltKItFCNvIsVwUFVCGUuCdqKTyY47APP+JOiyCH+U1EBM5cMrCEd8
KNDpVwjsY4bCEzu0zmZ9XQsNEjg+eqcm8AKwaYDIJfkgO48FvLrJuhjN+3VhmfmDGCqrTBAwQiB1
USiIkTI5SaGpDidI8qwAQks4O2E57IaLY3xEtvq289c4tWvZOX0sckCJuFwNF6a91taQ4ZTCkex6
pAbXcocpBnxoxsvnhCT7tuyJbxYOpl42fnEiLWMSAOBT/KFJ9FdSuOEum6X6Z8NNV7CfyBuvdO5L
iObYSqNpBbYEqoLryOnkH374AXiGiKpmpTa4i54QJ312RwBGFytBDnkDTaeqWIpe089utmHgn/4O
x2q4VVDti79tfKg9sqOCQ0B7H43nRXMOKdSXltSfIn0G4Z3kyyjMEAaZzEqMSEBjMqWg1egX9v2y
OcyE1YOa4tOQ20MTQkaZB59my/H1x6uiuF/jgV0ORmjJZNvDyiDDH/rP2oRnhFfllPuOtsDO27Iq
YXmiob/6gfdFNtsI41BUmFd4xL12h9ypXMjjEtT9+Ap/H4lymvH4cOIHC1LOevMuZ3JcMoLuAKMC
1ciwJ8VepX5A33Qy4a+VvSRacqBUHr6crhKUz3vkMc1/MfJgCk1XFtLyJJxY+NrGbWEcfBF6uxOD
TXxRIxLCKtfM2pstZisKygY+4kx1JXxDaL/2vec5MRN3t41hauom9evtzinUF97kNet4hT1AQa/E
NkGvBALtI6r3fxARyAURWRB1L9de5sX1z1vywSzoOZXZU5Dt3tx+2zJJe+kal3TWb+yfkN5iLrt+
jh+zM0wah0R/QtujW/DeWI9Rcn6946DgbuRvXKuPIzpJS3YLJ2VWtLxx8+z6d0eNtxX5OfeFhKv7
H+pOHteNVz7XH/AFPseX2f+AJdKcCuZs8SRaSudKn+Md5K6/imhJQFAeOka8gRuep3jYdVr9l6Ht
dqpUXr7LsJZ+KP154Y28GTGWxIxvBVZprnxxHSMa4MwYgA33stxh3YtiPFs9KhkJJLyn8eU87n1p
9VG3lIfOvxSrY4/1lqZl6g3qx5r7HX8AqsBcui3eKvgbfez1tRjIK2SDP7XIBq1zEH8iuTRtVBRF
KuUXkyDzuAFoEkbsUWvY0ppSjhQlPutYBv6aJdH2ENzgWBUFpdk1yCs7fzBHWfrodyxmABvla/y+
ovZliiLDrTHCbsFQOM8LqA4Ws+OV5KfDG9Nca/GwqoMnT4ELpPSNGhkSkM7+fGaNFrge03YoBxFj
wADixxnIh393pHwDmdpS/bEwajWwuSrPN2mj3H82voSXEMGbStqcPsgktAwP+lzNZpJqBumbLeS0
+3Jc4MLq6tXhaJ2LVbNweewHFZ9BX/JvGuMvl+OHWoH3caQfcT0FmUNx6mfaKMp3CutnZZAVB+ff
GB+hL7FsgAEf5HbIIb1Houulz4Tq5VOihDod2csk8hXspq4R5RO3crhORWvL1NREk/UeZuEtT0gi
j4EWEt19Pkksag5zpjKzjyy7O8gqrM4A6VVI7gvITl8JvFX/eGk6dMLZgu5kSKJ83Kn8BifBgNEO
oaG0PpYxuLIO01GU5HPPRGuyc0dmy9jTee3omoCMy5BHOBtEqpt//IGNANXffOquAjLiLGl0jZ8I
n5E3p5RaivwUusJWx0HEHAgVhW6qHEVwsVLwl+TRQ6ts3+baU1T/fMLjBvsPds7n/eQM3GDakS7v
ibzEMdqvVjynrKngFPR5xddj3wSYftXkIJChwWppD7D3lycIF/6dgyyjC8v5V/y1GvmlWm/roXPs
eicV8RXv7sQ9Xzxcrdp3v6Io9+P2roSEpJumDJhTSts3VBZSFQus2sPMEtjaO91HznPQZFOVKLsM
63+S/oyxHLTm/GqyR2T8Vo1uLT7M1sr090hNDyySVNG1Nu1QCIKY1hswNr2kORR+KthXF3tdN1Nv
jXPqYGz3Z9PU9cz5gzAhmb7ZXnAnjQVINUx55RvEHwmIBcWj7BnnGvwq8k03JZB6yJL2BODoKcSU
PgBbNV/5UhAwNy6gUzHjFdohXjpakiFQDbQvmZcl8jKAWX388fXykTAcefjyoL9VxDXC9VPZQfxv
5oF4iwMppeSF2CpqE7quei2JmMQu6CUZhGZtfIFufNSWVF+I165DCVHqVEIT1ko+EdJqeDb74Ytt
sx+OyZHynYybWRfqHa5koumMNCCOSS6RadYM3+FqNHK2QsuEM+EiXaTQ0oxq4GfRFPMwM2S3PTKA
rp6ws4yoJj3TVt3gQjzLL5u4ksM8PUxnwTQNVcVn9AWmuMLvqbqpyi3LhhTyAzwthzCDtok6vwXg
qwX7UUHDGmo9KnG9L/Uz862+muwifu9auNrM+lPV8DWJfNkNm2yXTTFriLZk4BaOFTBAfabf8ChM
DSmLsTwpAEmDqKQ/yOXE3ZTqDhVjNhBSSUyqM/RJ3UZxWIaeB3rUTuvPbAhtKxjxd+KP3mjpvxPa
2YvOeg4HgRcDgcBM6YZBpGyJRREibu+su35BpYAA6w1odsUw1ewsXDUmXLZzoFNSV3pQm/JTfIEj
au46ScS7GRI+1DgHby9cmK8H17ZFAa5ttQIkkKrcpfqE/1aVa6toRskPMmjmP9jL15qc9wWVBFG1
1cKtcQWPb7AvoxmqiFslCU4vvb69PHskCX5NbB/enhKwxfk2rs1BioR38hMOYshHLT//dRbJs5K2
9XLrfY2+bMNkdr/joQxNU6z3EwmPSoWG6cw8Af7ze2V6kNaRZKd4HwN3jwhUecc1K9WV9pilZXX/
1vONJ3aph7rgMUa0EkZO3c+xZWqLG15AUVf+SOX/wbrvUU1Ezg/p+mi5Y2qbrGnr9CZ1/2mwp+tC
lOqHmTWfEnf5SNd1VUz6rk2jZKph1tKYfDDgD+fJDsnmfjLL+asgDIAV8iySbAhUQybtZIZjE2DD
QNVlW/BruYpA3PmpuOgsOLA6wrOdOcg6oQnDKV6M23iI873gpaaP+LDpknbIZUDWsO54kpTutLDL
/E263W/+KoGZGdIHBssvw21RXYEVQsqMAIwXVxlv6xvZsu44IjJINQZiFeq//OCansv5S+mZH8Lc
qHny9q6kZNGyhjtPKJpRZ1XSR/K8i3esGbObw8Fqphl64rapa6Gm2Pu8xDA1F9Ox7FPeig9kk63I
4rZwZ33w7YlIV7n74XeGw917JgGJVrbXM+qhQE1yiFztqtdfco2SDUWyZiiimiU/lHKnk1nP2jNS
kSvundl/6hSW7VtjL+eRItL/iJNxaJ6W+F7Eh6yomzbgoGN+LXYPtw0VT2a4EgGk3DPxAlEHKJJb
LUmDoRSIGBDR4j5UJ3FP6TRWNffWgl70TKnpXlLell0Za868d96cTNCk87w0LPqhvH1MJyr7a1sR
4BSZ7Ib2QOe47UvOMx0KT3NvhGqeLaWeiddCfQo+C+Tfe46McksRV8x36dzznBSa6ijIorqoymjW
FRIuEB7gaNNq+sM8gh7i3CTw/1oOpCDNfBiJbIuVxsqYlF9h1KWxsg1WawivfGqrL7k9CR60MamB
wgt0KtuNd6nvvr4bOFTlxb/iKld68tnHAFbTwjMZpz1x6+WtEd1J+IbN0OWFEmAU3CRHo5NUwy0m
fJZLBE+BYaQ4VqlVB1W85zkNi29+RmtTwLkqQYi7K8i+lmMIvr0oY5Xbp4wPZZ1vK5H3ONFzViR1
oxNBWDDYFUVkyPJyTS2/RUNP27iph6FRUvsdZzEYQUOyPs5x9v+gEw2XHmH4NPeU7+vleMNtsjxI
FKGGPebBHBvibn5lkRIQNc1xoghfkvyBrpBQZRQ0FqruoJF98cmQTdllguiyQykI5HENCudHPLIj
FqloD7Jsx+GrEEr0Oh4al6Rd2S0KLHLmb95CKJ13YbjDOlHsmaL9yTQnNwYZz6fj34pTaXKeDwxT
6aTrk3/0g6gNwUunx9oKdbyY6A0p/SKULG8fYkQpOqm6Pr/afjF+CiyaClyUZFTD3klBuzSf579b
bx3g1ZFumA2eZrceWDuRTpC5VzPNkfurQW6E/MbSNuU+CvVVVN7DPJK0H7YwaH2+Ys6uXiWtBa5W
B+TuV26Q4IL3LZRjVvrMK+5a1Xi2E9WLZHabNTvwOk2gEuCKOj97zEGfssz8Vs10Gzwi/gYAZDl4
dvWEt+8LQq/0schqJHqalspG+uQirhXEjQ3JfqLh4WLD9twmDtB7HF3yLGiTg5A+1mG1VpdtcD/C
l+KEdMYhbhpFu6I9qtg28e7mOx9Li9CmTtjcNSTnj2mKs9XLibZLvtid9g3v5iq1aet/1WOsrj7Q
i74BQvG/WUZhTIbCgkkyFKnLcJhhNMPoaDhlBBcdWZOTH/qxxNycYWDvXjnv5hO65aseDrwn+er9
hjq4T6ETMR5w7KtwJpBrhnaBO3l6C7VHnNKfnnb2DFJdW9qb32r0fQ+Hdm1SGZr/mOPCKbhgYEnk
Puzw8ob3pKhY++6gi7MlXpJsbxPYHMvhzrnt/V3693AnokPAjLpncVW4egu309lHl+ftucaVzlXi
rmspU3AJ2b7FjzBXO57fc0M4gCUGfiQGZeSt29frVgnqagG/62aq+3kY5bi5xS6Q3xm9+OdhsnbM
1ccQevFtIcthv6ZcWcLgP8jEUzOZLEgEXCLoIjDD+ED9ItvRZkogUInmlVABUsLOMjzNJqUpMk1p
M8orpGnV63aF1BaqJyhFcIsUEpSdI05GcC/gfBdNYk/HMfmf1twfKR0j6FuFGv7+jI4Iltpvh9oj
NQQRKtAGcZBV5j3rLS6eI77CrcN4Yn2YTlRhyB4YGPQq/2Nc6aoG42O28FKN7gag00jfkwC1GfdE
qzjXj17+XexbhAb6DDtpZEaHh1fT+DjIl/ZIxUsX2qhUmiSQFfss5whOQ9z1gEKa1dpmZ2L8zKPW
QMIcuenPzCqkFSeA9c+9nGzZFxHUefOrHAWPR8G8NHNrmPHzSV6UTw9L41QPPYUoV4pXmnmD3NIn
WM+9VVXX9fqTm7DsSmVZLGHTQAX8a0Y7huqncPhTx23D9n0VqqPHyd1L4V2MiUM3bQxsM8Uq3/jq
GqW6dCNLNDDi57WRnGc5l7NigwilTvmWm7LG1R0Qa2z5eCajQXwXNGm8r6JOlyJAHjiFH3ty7sJl
Gae/WEyjQBjLyo6Do2ZFfr547pGIR3jkJfvqx5GWopQlqicXFlS0fVhKL28kkyn8ZvRb/wVZ39hA
+STDhPjQycIDlcFm1GtM1t1zGGk5slouOfM8ZIyq77vCPlXAYJTpN5MXUXUVnilIsv8UljVhf+Q5
WEw95ih/EY5YvWZeGKXuHwAcvD4/UFrTYYtocOTmiQ5UkkC3aApVAcrGOjMS23TSsQwCZKsnJ0Al
n5+miuICtgs/jWpl+hfpkop7o6hksdB3bX5uz3LqNidkWEwjO1x6eYGRDx8lE+vFN13/WoWwHwJr
DbXJurFHnzcQyaF7KOW6Z7EWCwF1WI+MKmpa+uhC6jjAUo+QMLz2Te07uVlaUi0zUR0FQ/xfHge5
HXwZM/bLFpy8rZPOo/AZy+Q1TCKstZv7xfRr0+Vbmzl96mu1OCV/g7jPv8BndEAqCd9qWX5cp0B2
tjGHGQRjZ2bPaE4+RA7ZMLhzDSUmOayuq4OfuKm9mPc58bIPoyzFvre0WSSH7YMmkucO8yo5u8eh
IzrAQeTErh4y4LDWoGnh+ZYNqAaRLgalSwJT6cKZ7QDEd+75o7+nkjI0BgpmL8GodQVIoNaOjTA3
pRi09W9JgLar2tRj3s58BDLj/GFT49pvaOxqVdTejUZ4/4fuAuEU2XgIhA2rafnq70hlxmfzPmFu
BO0RYDPz5r8VItPGtW5+bYvXifCwGNL99KE9HrSYt1sC/6/GSfq3adPVYBH9AxnAiaZWbebrBVs/
DzsbXjGnE15ZQw/IkB94fbSgCiGBxcg8THnMsK5zqqOV4yaGBgwqMV+TVcr6tVg1riJcG6uqQtYQ
xBBt/ArjwDqqxWUiqbXxcHp93GjIBhVlo3HY7RhGrFcnRsgnQAd3u1bGlj8ATkrUlqxsyYaOHisE
WpfVujCDz7yIp1l5fnnG3Kjzut3OA0084eMa4JT/H9lKXnUHh1oaijecQHpAVaRSi7s2XblUaUN2
QVvHeb5eojhgzs1fjHOGImimObSR+14la9Y8hIxXAJWGPmd/AHdQUPw+Rx77zbrJRjzDsa8862K4
4acP9XXY96ybPA6qbO63cWIfClxItMM/2Uvpix5hRNEL6IdjtKQqqufXj9pyJNPDeIRh2n1xgKZL
527nHnCBNivtnZOmUHpuuVZzU89bQGYsoPRUuxRxO4RoHHBqjdTZwpr0puOXXic44X6CYOk8y79s
GcUw4j90V6Agd82dKx/ZEpIYXYnIQTtrB28jXj8hwkrRmCdpfVD9dqDt+Fy6krY94D/FkcRGMUWx
dMX6wV72hDyHFfGEF7ISZRCrPJqrbeAcTELUFj5YsQUkvqGF3jF1Ke2sU6M0TDtqhCNfsUJQ0xrC
lrJLDWpj3pmf0NMRhsVvg8pCauFOoE2tDuGeUjiPd+t2t6ydkEBtpQ3MUMixCoWJ0vGt7DWEaHx3
Kbp54HfWfiXxCo9TWlXvpiXOPb+7hmKn6isq63xSKJvQGpNcwfb/nDzJoiya2A+b3JbGmWolrlzS
Eira824NyE+E2IStjOTVi0ZodFGaFCjmhmviS9bOjD/5mGhuH1be2pBosg8pUCn/IUFcn+uUTb4P
uvqWfXcb1RCh80zjPWqYtJYxDu3CImR5HtpvrCRZ2O5/RhpNUw1C9+vBVsbDMbeMYlQCPt4uySHJ
z/uleXFulGHmRGqIlqi4XOwTrU2SR369GNAHARXGmCHhB7ojGZ7VMY0BWT/LYhMQEsft6jEIkRT6
WNrFzHGPIqGIENpOVv9IpqoPRM6sQj903ykfGX5W+HV/UoeVHeNPIo/RkbaI17MDgA78lINv9u/p
EZ769o8xIdBCS5hlk4phovTmjqEJoDUok3h0QhINkYiog6LwpPKuIAWit/IWhigsyTdh01/kO+4U
fqIdp0NkJ6PUh9ZzW8UxkerOLW2jNtUUhFOPeXV9Yj0w8uIPbZfDkhtyL9Wr3xNBKEjtLRV8yVWG
dGZWM1YNIG5mhj2D+GBB3aZ8O9nqQJ9D7GXDMX4N3WDJX0UNVGcZ1Uha7FYURChXX3YZTaFfI7iV
JZD232O6dRepyzeZ8Wbji9ps0Q7/13etNq2rFZI5QNLlRL3ahqmBu26UlFTP6azOTrcOSUF1XNBB
UQb6Et1HjttqMrgRf5fK8ksZi/zp1jRcuHEfzzluK0bOI48cguy3J4kZlN6HoG8lu+JDCVWqpIvn
q/khEtFoS49mOsk2bRvpFifDFovlhrmMJImTn37ObUlW9Gk3qnSxiAzNkDDJTnliG5gC+IABpIBg
/RUDEQNmCnJjwX92MZUnyxY36R+ZgDpUGV4QGFQJvdaSTEG/3gEOaihDibwtyGYfcFZQbJS6pUGR
AETLz7b7A5ySApKItlt65ACxSi8VMtbZde2MYEy72XgMHYrPs5Fgzj2yZ3AAlzW3y+lUIeX4iViU
XaiH3UPW4ftMWAEfEKQN47RBht30MWnJcSuajfQDK0I9Q5K2FK3Oqlcfe6PTZSITj/qIG1Ey6Izu
QOYkc0KAWopajc5efPPq3SjDcBbxvI1J3AxD0BcX4+UpFGHqnFamvyqneqBAJZYsL/xmkYUZWYcL
32ClcyDTOtAIpHqgb1xE3MymQ0sVPKxF9fTT1f6/PirqRQLQcj67IvcIuU/1ebN/SeFokMstTYFQ
bxRIYt3nmBsqnii2MFfa1gZM5deGh2cSicUfk6k8/yc991DTVk8Mbwf4wRyZrAEwVk4GlZ7V6qoD
3HBqw5kIj4RnAINXX633LASqCso1SWUWz+TTyP1ADsRK1aRuSIu/QceAK5yvlRVBL+aHdFXP4KNb
fcMUm8Nn9idlU11328M6Le/GPGEZFOJs18D24Q3NK3VBfKg5VykuIIUKvxjIWE4mLgbbaq+xi/s5
6hOdBKoyxbn9BwjWEzcfDnL7RIQQ/B0qqTiKFrZ+fqzbhdZyJ88x9ArfbcszNSVisU8SElnhsUZm
pKtVyR6wIK4m7qyFz4Vky5WJZoVBn988B+qGCoAAVpr/qcN829Zn5oZT/GKS298aCmg4QtHApTgO
KzP0b+V6PndjZ0dO56jPEjezxZpecHghxxiiwdt79Oextj001ip9VBDcTB9pGqJl2TTXTpAEfyuY
lq2/RIUa8kwSuWXnV5JcOmElxgjU/LVtPUm5+c48yyYUc0l9xWw5o7e4BdnRqN+K2Bx6QJqjRHJk
DlZ9iOteHRgEd2OfL55ywPrWle6l3geq41K7wBHpjN4rKVE/QjPkqOjLZsJGjv/Nd6NDWXZEhthn
i+fSR33G+qc7iagIQ99BLu7ePnk8IpOyzdkxxizS4n+osO5CVK128iF6fCswqGq0vf79QbO2FN0s
f5Jw0HjU3HjFWNh81mCTOd0XSgKQYtqBHkAcOeavh10UcUlRnack0+1xKVAJ5QKwUbr/OfjjJ0Y8
guh8L2Y8GyOkH6NABtaXJPL1rKNXzps11WbODjUlao5LySqr3kB0ZxM07u5qpusqm7Hs7E6wdrY8
TEwkq3dqbolHm2OoVnYQMmo/LIMMAdC/UaP9nWRGTzWhPkj6E368eiUl74938n1qn5Nh0fSHvdGZ
jJnbts4Yd76XuTEPYR7yV62PKiVkyVOiQ1YzdtLT+PI5ajkyVneQXrU8StrnfdG1sCQikNpOvyHR
US2NH6x11EtjYcF1azu9cYMiqMaaJmrkUVXLoV4qCEjQtBIHffFVFccNrJMt/EqL60COzrn7Pf59
yR7eu5k+MhbzX6sOOUjDhMZdPnuJsxOHkfktU6uvF+zCiS/K56K7Wx3bhpD/erKpXGC6ZetaZnYp
OVmMXimsizMHZG0O4TdXf3T7nPkOjuPdzmLGFgwv3n6I7JEENphkw2ME6J2buIvKuhPqnq9F957w
vkqNN2Z3mVCXisLvbgOLfp900nerDMd+Zt8E7Usf0zueLetod2u3+6yRplHq1qTlIfX3Mxp7z1GW
wkB81UiiHgJPP8aS5vEjYjCAD9dAbGAi9tg4Mgb7Zbm1Jx+BgK9/YLoINt+zTbadFeqMOVABjfLR
i04W7zCTpBJkAbWUag0cgOF1xuGEj2ZX0iLXeJHeTPUI7vz8qnDZ4DgLS9R4BIVFImKD0Z38IdP5
q82YneISb82vT7na+MUI7ulqIRYRqmn0ZZSFiVwSaYhlJ/dohmdEIelc3qORyT5/Xam6f0i1S/DY
jq2eCIxWn45UzO3dUq+JXEgdLI118/XX0C0a9NZMCuu8RbsP1wvIsgBBr21gMRFvcNyPfemjEl4t
4GvE8Hqc7T6sqBspOX+By4qie5Nq8lvXwGRDE3YrQdYI1qq9Ke4taJlxRQnF+zIEZ8FDgxx6Sl2f
vU+ZDu6dNEMDNdrZwmawSqLUFTpRLLkuKOH4khxQIumlfYR+OCtLKKlCQOD4R7aiR+xeWWD4+hnm
w4YslgeE5eayqU8qvsN6PChLjkf+jw/UDY6NuYrGcqODmdaWv/uCmtKVGvXpjf2gGQ4lnJHflHvY
CEi+I+ib25WGPZjriStfL/g2m8rhjBiIURbnFVmgmoYQyQuNs86kzpLgAMQghCryKuk5bi/eQX1R
4V08HD3FOGKQb+ODOUK/N3an66uYqbsFc6tKjn8h4mUk2vo4CuvgM9BwglrfjCPzAUtxO6+dIc8m
7Kd8iIkFDaviXn6hu/i37Z7AhfcrumChTh9C8ROV6XE/jkJOMdEWIQLn/Dkh7Z1esfwy9f0CPYnt
+8ytWv8TD2SgfeztxRTeT/FO1YVLS991jqsW4cb0WjdsSy/++jNgZE/R7zE7Vphf3JICWLw+ZZ55
fEa0iQR4oIwFRO56bfTNbu51KKs8C4wMliYUH0IFMsGUwG6BS1X0mqGyB98I1mltRQpiejU66Pgz
5LFatw2NbeTK4YcKg5YVRb8TDQZK3k8LBrQRnIwCSY2Qa5/qCMaFS1odjinq2rDUmEimWRw7Z/uR
9yUCVLmxIAusrWrJADMjyukVHcRj2umaxGx177jGZPgAqpM+U/zptXORgFQc36cAfw4ptzjW4agR
tAPzvDpALXlkyzmMhiy4bQayeTA5dSv2dvR1N2ztl4AZB8khfkhIS1dvaLfBzPOcIJoj+ANxV6X0
MeETWIpQNDgX66BwPAs4LM4HPRLin6PDegMLnfF5mKf2PcG8YiXxjCEpudwQ2TJXFQFWGRPSPClk
kOEF032tcfMzME7pSJ9iAgTh/T2P/ywmXX6fetqm8zpRZeFp2g4bVdEixbmlnbGzBEqs0Qpca2e6
Fjj54N5AIp6edAMWyhJrQUQQ6M3IldcldxR0VhkQxLmpl6dCZbhigWzdnBfFwPeouTfru9UWrIE3
2IuI+pLF3OUHwvIe8rLcVv8CKLJsGewhbW6h0B2PbaKWgnmWit6kWiVEiG6SlSsI4c264fTYEQij
rI0EwyVtivjok8R671MWRVK6gmrAuSOlu8uwTtImSUl9ThqpVHKqkK01xs1t2BzpLQO9atTnSNOV
mhrW1p0cNSWE58rXxQMNI7r9DNDb1k7l5n0iPPaLwOonNN+OOAzG5nM/e80mD6aHXrCqG3LbzKI+
PTJx/bFZ+1WYOMtiz0q9r6M+MeVtEcYJ1m1jHLUH+uBCQqOFeiYqoPVQtk63BlLYLr4DNfPs7C42
qpoiSTqwvsFWB8ttaVnGKHhUM7VWWae0QwCUqTjGxnMdV2sbvsaLWKVbq5Sl8k4NBtJz5UQG03dw
bLtlaE0XndLxVfGDbsu44AMs4cZNUgbEl747fQ71ktsFD6poJ3+CA632hi3byJcCeDIGNkBO7CkS
EbqIhMpZfNp/RtQwNAOJPoCT33Dncm09XxtiyYU9jTpbjRNRk/ss2/DBzfvYB+MLI08/IBm3nMOo
adyR3rTY4kCyVwSCUqHeqg3r6xLHALixg3f627hFXAO0f/TIavh518hbiZdpGu/huWHNQZTNgD1x
YXcCZ1VLhV4uZUovU1zsI82VV1k+4z/yImfHNqmOHcoCuH5CfQ2s6+q09EY70atd3y950e8XmGLE
B4Fpdukphnwel8Gzo1SXPXfj24O/HbLT+hy4xVRORuBb7mVDcSS27VbjKdvvClwEAvRSKO260luQ
IE76wrlSVpdTq4Xe+87no5/jFGxw7eRZ+VVSvNojRXmSfm0J1BHpGlG9B2eyWF+M8YAuPYzGpeqs
YJvNPnwGqGCfP735i5r/lBDTmr6YDNu+Up7PbuSmVjtwdqzAi6O3dJpkkZZBJr+qfDooXuDPWHxs
FJnIXJ2tLd74YZQFGuydLM/HlLTURqqjyi+/277Q4Ez8gtBuK5dBOSbGYiwjto4IFgLxgoM0jWr+
UEJi+Enk76vb96iFyS+by3w4EqPrYFUZST3oLWw28xpk+oOgetUpUv8WIQP0UeEgWaCZr/b/wm6P
BlL4fahPYP6LY1FJ1lfmJNu3OH41TyUZ+QorRyBQEY965G8p/2O+WOuLEJe4UhtkRPG3sDXjMIx8
3o/AWdMidshrBto1HJQV6pfJi2NncSYappITqYdt5nRRsMihll7l/ofZWcypVZcQF7eJ2vqSUsrU
81W07v2/6fsiiJ+7yBE59zTvDR1om6EgAew0ABL7NDDpnp5xFOm14VYIWlU7yfr3OD4ny2+DzbqE
uAtiKtibi1RhpAu4+6M640EsrWcw1LsA5tXKKifSJF5w0MVRsY7iriUTCdNkWBdmbhGMpEFMMlFc
vYTPuNFCsvMnpYqpP7b1oK2cOzCmD7KFo0OfprNA50uXPdTwFKuJ7fp1+qFYXYwUZ4bGQXUWxYHV
XhHgpAgCqCU6yJQNaV/Tn3DFRM0dzJvYpazwoSYiUacFL9AsNQ731EQCC8N3kjxEoAocW6qAsi3X
IM4LacIrbEEOP0zQLcF1d+7JnsEqtUbR3uEsVqY5Ub6fQotscHKrHvtFDEZKPoWX/JX+B1mG9lGv
w8eGSSZD7dlNwXMz53JKO58M7X7LEHDmZrP6l6vRfvzHWU9zHgdK2ESSQKhuoWlyWYqGyH8dd7mD
at39LGohkO2Zhh3k/S+IqyoaqJ9ws5m6BcPY2K+WTvmrRtCQorxvlIxjFItu2J6qYARZEJklEaNk
isKFZHvSyY1N+vBhzgGdiE6bFL0pdvlOOoZk0a/cBIueX+/UEh51RzNLAMtxD6OJyXLuOkwL1njg
iHPs+aYibyLAS9qNnbi+FGntbsdvV8OjMyk9v5RTkEx/GDzdVjxx3ypwCjYrXr9Cm3P3qVx8ZKvn
Bykpt5LBznoOvZoAH0qV3Bc+V8KP9VaMqD2J0b6m1mx8DuPhWoy6Q/cH72dJboSGzlzpvr/SrTjf
6WaK7RAQD/GGShVt04g4hzCjlNqZmrtN+CxdI3nbszHQDk8e9Akzwtgx1AzrM3LHNZmB8MBZ/ilr
+2FzfVXz+seKDDly7WAxzO758lqC1KkCXwlcQ2RYuWNbQnAUB8bC9bHBvU7PHgulZ//FTTYQQvgw
2pAJbOF8uD/QLgAQ+SD/X1/9vobvcgYcBkARERk0hLuQqH1t8srX13NlSheoTJvUH9j7T/we1P4o
Nrjgyu/GK63NflsjC85DhFJaQFsMraNREhbML57y8LHPZ8mYMB/NwWGicN/hA5fBrNDwMUO73zS8
MFxGOBbB0RrTglwF4A3xgyz0cltt6xXbvTzplkj23at5gLMugWUTems/Xl1j3AkVGCX6m2qk17hV
6x/JGDsTIBtGPOCcgYsD8jd7d5vOI55kCISCFle5jfO5+wAxY5NgwbpApyHBERx6rE5gv7PehncR
PZdAOFpjydJF2wbypc8CHREBf1WN2ji+Ksqj5rAGnhjtqe12n4Y7K8cDUyHEaHo2jmVLb1A8F3ij
yulOIyvOX9b7Xocr166Y9UxTCQPI+BFvewZ+LVu2wecloNqfABkPixnyIGqNP/Oh+e7MHzxdkaCW
urp62i2PqRL8iVFwHUbt4NioXpke+NlyWk3ThG7W9gqs4Q3GFbHFQbSlB36zwX6wG9s7+Kl0+0GW
F3vKIrynCADlmM19gHeGfmxp6a3Qh4Y8c4EbTPK6NyQgdJHuDKA7j3SymfP02Y0MAZS+gg5/acHt
3blPATebXVeKQW9Gf2ruGMqfuSMdxQyrxJMtmQYpY1X6Mak8ds9QP2DnxBRjdkaJNdc5bGfTgTNP
dlQyYpHimc06KmKWCNK3vXXK9DcxTcsiXn93LMWqrg/4R6iQq/tEm4MqKZhdzkNVe/AxTTNl+YN9
iPsUgq7pCRO6d2+rqH38fxhSCnxMT4xiRPt8a4r3CRdFoM4ZbEl2Jtp0XQ9lYSjQvBPLERa4Mvfg
65JOPcjDjNPoqhfhwB2Q86s/1wC9O0zUeN/1V/WMpqp68++TKVfi4c8Y4knSv5JGijqFfbEu5h3j
Sw7Ks3O13S2xPTbk2aFFaiBXQvPuI56AOethA8InAIIDKBUcpos1iKq7at80JF+9/E+f6UwaHv44
aaFMzUDXw7DqKpIfMoqbT27azkmnQ9DQItVZ07d56A7sHI+KFhE/LZrRbv2QmzZxMTQM7LiDIK+K
bh0eD46wxUUQZiR1IUil6RGEVo9zO1Td1RuqSBomPTzHrSkDjbHcu+L9dEN9I4AwTAiTdXWwykyf
SMFydNh1UuLxbSZmnaUyWa4jqnmm/6Oa4sgD3OhFiHNC3MogjsjoLXdkyP7/QVEN4wjClllOzDOo
iLuNKPKN1bC4/PaiO+19OkGyRHrEJniy5cb16aSE1NTzWlwJPitjlNVvYAWy7krrH6QrvYt4+kEO
oAK1Fpiv1jvUt6kRFR30AIJD/LtidogXglNF+yz8BegzidrPwKDeexEvFmBHFOW9DegjRPq3zEVa
kBsKunTEJPduLiilKhsD273NwT0dgN2U50obSKYn1eWBSeAakQkBFHEbpL/uq5IuWnlqL3mk9qxb
cULSGf5DUrRchtDb253PeHDff1yU4kDmLaXafxj6B9KBrwOBKCs7xZjXyzvk8qrlphsvNLAjuqrQ
BvEBeu+O+r8S/p8ejVNwZAClr0hHXJsS4KH1CuLxOkoLRwtQbbrNSB+PjXihA8mEBlonKig8Jv1T
pHLyXjm17XEMqyCizEzzd3B0KuN0WA3WsVHbzPSKwqgg4qYbNTI4V5vtM6Cku8BoSR4Jp7LztCEl
SS70ix3jYa7ywr2mJ+4azCerA2MGM3Rn9OjfSlxlAr2lWzgiYxYRYdoKxHQRxqVeVU2a6ErUzZ4F
g2gVTT3qibHEezUKvZhNwKCHGrumzCbnriTsfnFV1ZxS0Fcz4zfiYfEzW/vdf9djrF82KRR2v7ae
ii2VCy5StfdboFzg5ioNYKbOSd1DOyZ8RxRlPVTI8+CFlPGwj+rBfvE+Msj0l3VdR8Yh3VVNLi2H
3qWBERUOtnz9DywkGg4NEsXY/H4hr27vAueUfrgNzZ1fmJY0bAkBM5oZeR+bnLu20Cy3MaoEfTGZ
4lpbQW48gJX2NaAOvKqx2fsJWB8jZZbUR0Cxgz6bfsSD1W+c5rh/R8Yn7ARcZ94JVkaCJa61eQOw
CjeAKZ+rjnRtq7GGskfC+nI1U6Ed5yJjrHTDF5zjHG0MKzcPEKEBoUrFiqcAGAUq2m0T4arAINfV
Xa4I2vWz10vDFvI+aQeaD7S2Wh27N+pRyxFIOGChjGisWnlZ6ZMuNrpg1XNN9Qz7mli2iOZ0wU0Y
SJy6GirTo0PeKMnjHljTHRHmQw4asIqanXvqZuDMJfmtMYXZcFL8bxp2x1TOoYaqbYlDMgdvyPJZ
EedqoKjSudbh7/UdWhpb3FhFoiARnz+TMRp7/N3wU2ovQ4Ek17r/i2rST52pppz3wlMMA5s64JrA
PsHKI810qY2gHAEojpczzq54IP9S+rnSkvx9My46Dft2oqnjKvVEHjrvroZmBgIJU9hSaDAFhKo7
B1Ckjyg/xG4jDaUv1+FtqV++sbzVX624h3V7qg/eqcvyXUvxn/ITlQ0i7k5GsCVjNu9o9tWwOs8d
cckxeCQ03NkUPGNMEt4jy/WnRdNmVqENQISm6OGTMsaDnXcbGsaPn3lA86I03jHIrj2UbWq29tan
gZiCMth2PhD67BFvHB90vM7PQtYA/zS8srvN9I2Gqygdqol7483Kmap+Mm0eJfnKQyEAbTjIpmsy
z855iGxV0icb98l98yPTC57U0vYYbTxaVbrWawYrd4pKbMxKYV2jLMegFOujo1W6RwLNJFEIb6u0
3qvvvvfmf3tFj/DgDOoLO29bQhwPONBWicSeqhYFX9/fprJl1a69WYPs8q+I9Yzhc0BF6DOL4dZ+
EJK7Dl50WwPiwGaScpZMSSulLU2QrG6q6yzuL0LE475WggeLBwcJXeCGODNyAF8WVLn9oDhIDXSA
CT5cvoG7qsGowRF6i02yYVXmPKvhyG42zZxP/AuEulKp0vd8ltbPxSeC0z/wF0/3TBdgdWDzd3EY
4k+FCM1o/adMEtNlTJ0SD2lPk4qzg/V9uVNWRpkcEYyUNLS3H2rQnX6GMNLC79fQLmDDF9jWpO/i
FT/4xjAtB2rkha/R6GVaXNgtvkXtPbGYjKl1a4y7dMBuQTynsDo/l0LvXiUP6CNpTYXQKTQoa9YS
pJxlafzN934haFs+wU/MDBzZdckEpLV1IeVjioSSOzkIgOVw8ydT76SvMV5atirBSbhuwe4gpsiE
KMLrNT3+ddkHSUyu/IJeiwLcQVx5WwOQW8DrNkTBwF4ielFekQVCtTiRRYP0ka9pRZ7WKfPkNMst
30hVN1TLyoWr81SIQ+AVBO+8ocA3Rik/9AqtbYdosflYLeJE57OWO3iKz+YRqg77Vr+VCOQZPtaH
d1jdEuI5DxdVdqbXkK5CYT8PXP8rpo8KL7nQGomyYpzSTnAw5ztJCvv54ZlnAwxoP04jyATLwkSS
BDymSvDO5Hl0sxnrrLR9u45UB5Wra7j7ezy4KDdo0RPE8u6bb8xSFgkAHA/EPqLRgga0Nt8kvAzZ
i/4WW6yPR+48HCG8IYbPo8F8HqBjmCP6Zq+xNk8u1K3zMmU3D3U6PPO0WrTUCj/zW06yA/kYOR/v
82t1jSOuUo1n4Ly6F5xAO212XAAhkMOziTlC6Uyt2IGWMjLQ1afJK6AI/fvHvrkceJoDOYjkTYUl
20n7/pEQMPRkO2vfeTaslAgInRiEjqEeQQLyjBzO0ArZs9w+hToMz/LdHADm0zpCqqoQMFyqMYco
KsuW+T8Ec50iKS8ehEQnjSBR/kVNoSYuH9GBYGmbJs24TAH64mOPbSFfBlVPqapnmRcPnik/CC5P
Eh+F6ebH3oHRFFB4rRu5lnvT/ub49tZwfYXvo01Jxm1XHpsc4akHd3VOdRE6NqX6gw8hc7xvip9Q
06j3KJqgvz7evynu2I+oKhug3US4SvIaCjZVG2VEcoCbfqV5e4sCQyYOnWe8FmM/aThQKJeVguIp
vxqQVR2Ii00PUj2Q7oHYwB5N12ZltFEuESnJF5VXYT1Asgh4c+RhXPUO3zZOvWX9ktwRL84ju/e/
KclwqC3LGV8pgjkfSPiqSByqPym8A3alWzGlTvC+TBOAG8kmm1fYKMpjzJc6/6CD63ocR+L5DwtD
akY1tPFg+EbaaBSBmxFo75xy02gZhORrcS2QtOpr2HwJMQMaQNjkj1hcg7r3/n7Tr8vqM4IGSS9q
6PYEguL0MkQgwkFlIJpOKklIHRjPY7+MfxFqAAd++6f681mPQW1GxolFfJ21PuT8IvCXps1z6OaF
eAqaxUnJCeR5m//G2SY7JW1g5Y6l7w1zR1OwSjSnAgFY5dP1Ka7j+79ymROpjpb9ql+HjcSCW7tY
b+RNh75kEUd+hc6CkERYY9qsKahEM6iR8BbWhfuOHoxI0iS1nq8aQCUPkgbMNmrQj19FS45Cqfp6
jdWTx7mszKwlwUgJqKSMB13iTjZ5/zcoSGphPZxvcBHZOM88BVYzukWf87as4KoHR1c59nG9rXps
G51A+rmvT6iBjkcu9dctIi6dZlTC06K1xhKpqcqKbYdEFDLHoMGIiDnhka1gk31Q8wU/4hhQ6i+n
eODd+IXKnrkG1mc+BvXfIzCp0qn6CmmaLqTqvHI51i3LjlKV/owLhH44k0slFXYRxZPEydiEAH+L
i+5KaSyxObqZtclrwaQJcI0OBi0+MTzFiBd7O7Do1ip4GBHNq7z7rQ1lDWZ9eU49OunGfW5iYq/X
RYwkg/iAA/fLGjW78efxxyWYJexSwQXtM1tz4fQOIsZFyRBNWwmNTDM1af14Rr5oc9San0ufB5tc
Dvfs0aHDUZDaXLC1eGjBIHIN81V8x0X8LMmutunTJda/uT4odKi5y52yEOCyGUyDcdOu5p/F72na
U+401XxwRSsS3G6JOskjkg3GoMGRmQYcGjQaBdJafe/8FIrl5n2WH/5no7lby7f78PFuoz0yFp/M
LkldoOW++oXyizp5naQWDYxf13USXbn0y2QsrKTvyXjlGZ6JCap91HvKkWPWIE1AcRcEyZSkNGdP
vZxMptlXxlE2cmeyA4kB9hod+UndkdQSMhRHtenlqP3+x91cNMQpUSdXS/jBuiFCokVTBeBBiBCt
E7fzuWbPPh96z5dhNI9mw2bLdjgko4aTaFbROgWRl1ERuM5ZnASISIzrGNqbw/OEbSNTsLTbFTzs
WFmdF0mMfoYkTD5jVK5BaxebXlAAxAMsyeGw9v7WWOh0yxdI/nxuhU3Nf4MR3sRCLNQw8UAm2bm8
Pd72Y7d8op87e2IMOWmxAjuUqDGO1Oy/xcNJi02XIZpwgZfoxd/bwDW8mN6LfMl6OjBMV3jNS4Yr
+YtEVHE2xqeB95ZReZcq/TPV4d5/o78iZryL1xAwg9bxSX7BnLEEgfGY26pFPKKYFSIADyMDwz3e
NwH6GwcZM0WStrwtBTCauewueyyiLlk082PmhHg+RQuJZ+Lh9YSycQIn8GuM5e3zTQrU59Yk+du9
i4tw/2edE4JVqNqIGrTKvlXZKSR1B/bNk3RprVAACxt8l4GPXSasdYTllHafyBhD4+3IdH3/n+be
yqQ4uc+DE65kQVDHko97DZuaexOEkx0Wr3zYcWBtIi7DgQ3YtJ6ONiEIQZAE3MGZKm6uC3ssDyZt
ULUd9gEcZv3ZAZmhdSBQlOqrrNMlHbbC1tYfcvMQ8KTivcNVofhwcAhF8vM43rBx1Hv7ByCxAnm5
EEYHcp16tZ94mCv9dcnX9EdH0+L9+bFyfy87J5jvn5WXKVsvbjdnDMsF7RG3O3SlKhHqnDgsf70+
+cYBElZ/KBwno3+zQ8itlFNKelxPKhpYCU0GiTODpqsLoNQeRnme//iZ1wugZx7/txnuFONK9ewq
BHHJ8So+G5wc9tm7uFckANmYHtVAn9sTZC8RTLvtAbyxUR08gPOm6G4XTEGrQtwBVjJRwlq8hlAA
6UM2ivWu8mC7g8fVL3/d6fycLxXxxwSkec+gxwIDSHLWdxMdX7FNSZ3AE3a3nURC82ftqwHen24E
5srI18I1KlS2fyHWwMDa2OkvmIkebglF6kZC9GTM8W806LB+jDxDJ+GurBHSuUTKDX1iapp4TLJ0
P1S0Y57NBi6IJVeJYpBnjVg5vxqsy/AnSCtTFCZo8ZWnqiOkTjPk8zxNI8wV8eeysw55pk46scEg
6uxIk55CWwzDDS/Yg5eRIgEhe389JSKqXsr9VsuHgKP2HqAvg1iEnnXfhLOJC0myrIiMP4rLdf4U
E7Wt9ZAJ5QUWLwb5ANSHDmVphqWmXMLM3Oy4xsAuRyzsduDfEYy8TFmaNIDvhN593hBFY0UO1Hka
ASiDISWSrhjWkijGeAvNwi17zeWMihKH7QZkpniNSuHrPCmtsFNRW7D7VTraD1baxeit693e3c+i
n0iBckenIMhfqDkNpOXPaXUD1k8U6cXEDHCOHl7O8P4Lnsv04remERvUsJ5PdBwlM0t9peTnLbk1
tYspDPrcaD/72SYNca/UUZ3UcIiwgMbYD/w596vGUjFaV8amh6tfYuDjKdhwBBFoxwWy4QBXthws
IHLVi67+nEBieAY9NSMAGeqwefLYSGfbunOXL98a8AyKa2EKsdyLq6WSX7ElOSv3m2uZ7Q03Mzxj
U321Idk1Eb2jI0LzjSB2BIKi4UR8Ups1PRv1szsDYW6hx/gTb0K/qZMlt49UZTAp/dK+oXDgUxwX
S3pdNIQnMc0OVyMvuBbrP16LDOt3aCY/J1OiaIm7aiE6owNzAqdwCt0vvzIA0VeB5sTagWuiuqZg
ZtM56wQZCfKOJK25J93HIGesETcIJUmphjk075CqXOCWY/8UGqIWoATYwqVlQSV85+r6pkxp+op2
9LJ77cjnvNh1KFdUCtmfbGAfDGgO/Yfl0TJdLPJHonW80fZdfePWBL2cC3W+2yy2LnKAGKfv3v0V
QcRYlyHmu0SkibzRyHafAcELhiNRmEB7tChesDJcTRzm5KgjvBW3B3RCHfXErI5Qqlz68BPl+Gbq
NSGulohLBAmo3Ij2gU8g+gXCM+0orkubSOh1RPS/2NOe6Hef6AaYQP8EmgHd/YlqmOeXpukdWbuX
F4i0fKxqHkAZgtsf2cy9ovWEKUX5/lrJjv9rEybt3+JNUw3d7yrEgS2HRgsVzeCBuA26Y+PZw9Bq
NHVmvtKMHLfB029rV8teFFl5+Im5R1aPcHH02/aAMXlLhU0x509R6Y6ML+Z4XhvMxfLdQXRKj7ag
54WbmWsWxHESmFEq4nPwMeIgAZJmpI2tOAMfOfZjTZxmiUIS6yvkrZfE//tdK2YrcXAl+nY0jx7a
JQn5GsVJW3KntZ3QLB61OV/JCXS2ZeJ04W4JwSTDeH6Bh45shh6z8YbR8I+gqTWvGTvYc+idoEz/
D5uA0r7zC3E0wDzOLYu0jzinFTynMsQW/o8/EHn33d1RUXENF3r1rTRcMkZNgNM2hRDGErYih2u3
1gYpO9WwewrBi5wsYNAdJPYyLjX+wRWuuR6+6ta0cJGxBPjw3wbW4OVku/tEEDSRU29P8wRpZq1U
FnNvZbLxGJbWGJFJLdoAG5HsuqGdRYW8n6caALzZMbLrgCGoMmk7JRhRyIF5KPl5ehC3FrEPFY8v
NNFyqoCuEtvWFN+cKObjUP/+iSqG2Q4ENIDaFxaawbNL638JjwAsaJJSKqIN8NvlFHMzCLZb/zIv
/DcRqkJHh6LVQv6D6Wy9StOmYuHZe/4NjSwWRcv+ilGG3wSI3NN/VWUa2GDy+edGGu05QPgbj4FT
1UUCBJW6dpgiq6DyPxXRlr8CIbmH3C68/p/ljdwW/3qt6D7/Z3JxbFEqhGj6L27/ugXgJ4SQ2uba
W4afaDlOLMJPBx2jamKEgCYDia0AYos8u/ieXuLXowZEErRsiz90Sc7ARnGjRcQQ0bOhUkwCKlUd
KBeXB6bwJsVd4aQUKkk8X6fd0eCkUXa4wLPrwUw6x11UqMuYHI6eXMkpAYCnq9EKdkPUKsbSz3+M
xCUJmb1PT4+NeQuRSERVN/dJbSX+cyVfXUuzf/9cNOrwE0Jme7riPygAJTWeoqelLMJFQIuug6eq
ilkA8U+y18rzsmw0SRYC+LjOjmhGAbk9e636QiBUCGgz6ztJ4XtAPyKyfHcibpHZDfOSgWO254Df
OqM679mmQCPSA5rxmibn0RlHmF1Hw5e6V+p+YAqCQhIav8ABGH9JSOenZiCXyP5K2XokeBcXpAq/
sGTDjTuKdLxOwBEy4B1dKItqIhyFBKkBS2WdbisxRXp/VRke3lNxZdaehdxBD3JIm/Iv6r/VoXOv
hF3bdjmxZ+eJd6pyJ4OUa6TAt2KO0T6YP3wdHejDtbw1L5pbTKbzBlYp/Zda82r7bPW9soAnVdd0
ACAHAthf+ESmh0oe1mtGFRKZOgD42C8BpeOIg7IaiuIQIZK/AFG9dlcyxR4iTMwZGcSh5pQDIvP6
8bFa9qJNmqQM6vYKruUrR7lRBgRKPLe9zuJdtd4CEme69nOPDnvZA+atofQyQgQ0W91pby2VwaS/
xQ7214mFz0rJ5yYa1o7NJQmXQucHdmaDaaEo/dXp+s13FaKRTS37VpmhVY3xz8MNABhbNPHJR1Ky
k4B/L3HKd7TUPfpNNJyeK+NtZptlJybskh8i+qDcXau6FUXM0cmuMo0Bd8yV7iwYUxijXDGLiID8
XeBhn5laKFiiofA1BsMXRWeIOpteLRW6+Jm3n4VycjvT2uli16R7rNFM0KsbgBLeVK8EB87EBsvl
mzI9B9q81D/0A0gvwSFsGgLH4PhNIx7sjkvZiGMG/7KDMLiY6n+9rlmxD1fz/4XtZAaD7uA83QMw
DDCo7BfoAGckp/EnVrpuusg/nvupIBXvT2CczAp4HnT77U1R6OD7be4xv5uS/FNmCPHqhiMMHq/r
kFAe5zLrOOxWRpkMfJQ6nCcRrgSLK2mcw2jMRSzYa8sdO7CEuP3GvnPIHCqFwFS7Qc9GzMZECuw0
RhqJnNbRckQQnldB0bAJkCRYBuSra8n/gxRMjwT3VF9AOkixXj5GKV5iTooYyzPNlRLnZMYSyuRg
i38GaeDOAJ6RalJoUy/NWMgk+0JuYobDp97u784P2vpq+KCCAE6YoKYNf/1x51t6HCemVvzNv5Ec
rnVasLRlAIeHBEBAe8lMblo3dSCR+icP4RpwijujxKpyQnkEloQshGkDLKGFBJZAo0Ezo7k/17Fg
x8rG5xccYhh8TCzdiaZXd1pF6FIhZ35QbOIzq1+bs98FJXoelgROJuS9LChmjrZa9V5zN9fm0RMk
ArLvk9JgaplLaND35f7lHixw1I4S+e88JJL3uphHuO63raREZYtG5+HREwCznyK1IfwzcUQsa9az
HpjFCc1yaOkZ6JWqCfiUyRcdFaTCtPIc23+AVsqxiypI+QiMyNj6oNWcI3TUeibnqiB8Q7ukJkUv
ZRSmX3bkEleDSJxriXKuWCJo+0lES1mvhhIEwBpPTPA4IPgDtYseL26dmPTF9GrA82q8saLN+N3L
gaVT6m1jjldBeybuV9ukC0WkkinqaGXYGvtsME44mtJ2M/Y8rgDSuUEWZETsl7cUe54XlE84QOxS
bx3F51tSUY0aFy4pfT1o0SpOvvcMT6PMXfv5s0dG1UfTLil5Ysmggp+5C/M5lySUt/PB4S4PdNUM
gsFCoNdkrabS9aRxPBbubITnjInQktYFvqlV3R2bMseWRUivFYAY9UrHo1YkstvrzCM9Vc3f2aot
/MtK1E7zAgPtZj5ckfeFt0ESM3BYhrA8ZXk9tUL3HMrZnKKUzI/iJfKUoQk9kTBuz08jVOJMxkC8
6CEOPHf6FVe3NB2XMF9n7L3vgLxwSiN1nGegktewPwAv42XfX0N/eIR0EpfnpyP+RT0xns4SQn6J
q3/hTF5CVn3Z2qT2fBPWfwYMwLBXWh9ZTRNPBJQbK8J6Y8NDe85nQG9fauw+4UMm553P6d0ocIzV
3MEQ+h3YtAb7RDMpKsMC0wYS5J1fZtfVA2uOFb3VNvwrbeMNBTgjwlwfeas6l4au1rdyKEYox+pm
X5XDFZ+vEcfdPBuVIrScbplVbRGTt5BKDZfCRxZJdks9YEJU2+uuFF0G7IlE0PgBYZacyIq1Dn8u
8nU3kkeRqz1dBQ7CYkGnAyf2bb4X44Jbw0mkgms3zuDF8lQjlq4hS4gJEU+u/rKYLAT1xemTqmlv
tftanNxdcMgXyFfWRvzfAbCtMGHdhOZ40DlLA2bu5brK1tcJx2TGIUhgQFyA7L/UeNEc5iWAIcwa
QnmZAsSuOt69or6feoo5hFixv3o/GAdxYRwwXu++NskTmHjYAq8B+jHztzq0EnKFBHSX1ftgpXN7
62rAp4X6XHQyDM0tTfhMzdWCvflx4dakRbvCTi+NN6JIysA0y64kGnGrk2iJVGjbc3gGatL8P6kZ
nzAXYR/46pcEyq3qEF0N3ThU6p8xDCpSyO9AQdoSiWa43FXoW4pmPfdya1GkA/fUqcUQW6Iq3uy/
qvy5YG7KbFM5/DzO+9nJYjDzPI0JaRTsrc2JiUTTqAJzQxIrifEwvAJ39SCCWQq1kVUPa5mVoHbA
eGwo/zWm58XbyX/mTddYmsvx4/xe9VEy674EL5yF6kqYc+DHTr4P/6Cz2w31g7oXP3dAJmyv4yyb
nlaCaIZs7gkJ/VYcLTCJ1eKKS9lLglehRYm6TwtvnrQp0LUjBjesxi0zQUm6EuZo+NIuvuKv+ncU
0nc8ppn8i8X94aViC1T2EkrSEdbXNdSqAfUZ4PsYxpxa4qDVdYD0zEyFE3TKpKfEik1W8X7gyQFz
votuN5Y8AwiA3Qrnlq6sCz9nK2ZKg7KnKIy7L7cVolCFxqybPi5DXCXBitvF6qSvZUCu+cLu+yv8
vk8vZBe+XTlAuYuumnDIfhNIob5BZEB8x99kkHICcHEn9EPSouOhrYWs0JfPRESNE4gb5Z26+ki5
rJ5TmmvZU23JRHoP204hNDl9tTL50RyxMv2JYvit5W6MXrqL/eABbaUaW2zSQTMv+k2ZhdnI3/hR
4kOuAimSPW7vTqjDRgOq3X2zu5a7tfzqLpnm17s1zkgi/taDepnbl+xY8Mxa1jVCv6L2kAFCzYBC
ElOk+2iu5H6ZeZxdFfKl1QLi+e024T+1x4U4pOROnNOF++/3A6ZKzH2a2ojIK1dZmUhjdfIHHLGD
3NpkI11HSB4OhlKus1EkOiWXeiv6mw9EOsbrltMEVDYwe4YTtcINaXJCgjgHYQUnu89GuE/e2U9t
h0vIbpmolTBpCEwWPgeAxLiGpOhlLqJHbkbeQMo6uNnclWc3Na2D3a4BfspGR5pLkwzaJwFoaZu7
VtkKB0BTvNhoZ/PdFgDS8JECDTc/wTk3p0UOd+V+hqFUywAEyz9yn2SfqYx9gV01YVm2L/LCY/Zo
5OoFclifW0DqWhZt0/Sp1jBSHRB1TfVaO7EdhzoO7MUQMgFzMHW6DQoQUmWryHEbX9nCB5Z+XZGW
gGN5m6I9XFDqUxvCI9Mpx0SlTjnDNTfQFG23w4cvu9IdJqkd9Ol+GNNbRmjQNgIqF+UVT7FFY0hQ
alyRADQXAGCe2KC3dxW3r1YOFgQJCDIAkuDspMeaiQ+iOv45BmGN90oR43wbtFHcyCsHHKjikoUg
oO4N4UV9pAzITjL9LhhmsuxKXcrEUVmngDAIsB6NeAAp4uNUdf1L373BMzvwOeF6L7c5SrYl1uXY
Da/YpoZMxhqCgRhdsaeW60R6N/vQFyvJ6kEwq2//VR4mMP2BI5CRxUahPbPvRWwx8lAuB3U6BaPZ
OvGBkWeXvbNp8ycM6VetdzoR/9gkh61WJk2l4+i3ePUGRGEJ2jq04ze+vGtQht9BZ9012HGythMZ
A1pf887RR4BEtPULf8nnGFcwfmUkj5WiNPaSbvZ2ncJI1e1/Z1itomHAlZbaWttiqPIQHRnYCgJ0
PFuLdMAZNIUJqEVsNW6BOGeeaGEb84N3FQ6k45Wa3Xnn6jSinGK8oh9OEWX25gcXEn7u8J/3abb9
K+LZmSP2AMox03Rjs6fkuO/cyGbde2uCpw0h2N6VLrHm9XXnBq4qyA93P8iv9ueK1BXYffqkFWuS
YhhLg5zxXp7DCsNaFX4i06Q5hIJueZ7t815zIdYxehfBI8OZs8MD7g9kjoxx3vFfkTnc9coV6aQj
I78+aJeM7BQZpGq/M3EF9tP07J2ryoL9F8Y2V9x920Jmza0E3esBBx8HC/bi5AQXQfH57AWzWkee
+6xf6Ljl95OL29ZSr4owknwqaXxMVccnvtpxZ54TbRgl65RwZuqxatL8Ntln3rU0hrKfgcw1Tu0m
DFOD0e3ckI+1WKVwpVij3KCkBbhyD4PA0P/sMohAT0jE6USjiSlO605aTJ8gqR+n4UWrz4n0osDl
1tRvin/sHq9TghKTnO156eUB0Cy1Zfg/e58A7YbQmODp6fikJhVbU6XitPAwZZvDaGCiKVE6sckN
8sQTT9tDMIAMXIrWy4y7nnO/dpyFYwdtRzIL0kz7hLCkivVODeIY31Kr3IQlzE5ms4N0biYZITfm
FhGwyPtGbYlFNKqCxfDittCe1ZboHwZF/zu/CVGdS0gJnKwTwtf7SzWhFJcGgvkJTjVq3E65w/A0
k93XGLf7mzS/e7OGMEd3fbe8OkWaR+6OH8uRAvF8IfoG+kFsisyTfZ6mIrwI24EkfFe2CG2ux45d
yH5fyLV39qZpSWw8dBfD0EJTjdi7zBf59UHkok/ZgFrR10dE4PwGZIi1fMXll6JtLg/yqZmEsqyA
urPR/0bq4/uUNVVGwIWi9qQNfHYBxrsTcpZ+WxCrmyEF7s67/qYO0mA+CoprUXBFWnOVcgF1Kv7e
l+9MdHPQihzB505eKSeaHX7jTRHviVPmuD+dkkk0QwjAqEWZ5ja1Eq0l4sSYTNmcrYkYQ9PGSuQC
Cpr2jcoUIaRTesCp/A80YObj4rbYtHB8kg8HMZRyDgfPn1uFn1TaWJmL4p/HpotcVe6i6RsVooTU
HO7yp+HtGx3UearsewKUDQwZOWyRhY+r2WigJ4SqruQYX/x6HE8x0spsovG7dBZtRP8+UPW/d0yk
UXsvpWZS+T4jQ85g5YOSl2tgGGqphCoLk8A2/1U1Z61PwCDRblARwewJTL1KUhbwDPuUJaaIB2SF
ao+5H5B+SXTgeNOZjkpSVjwB0UT7uZQhs8T9mp8PIjeg/T3KDZn3SyD2sNnKqtjEmWLSWdygNENC
IKWH7Z+wd2f6DsNEmKidUMcEIpI4g73TrbMgGfcdek5FbPpzplO8CZBEhknqnuu1IYXE/O0ddkYx
GycB+/3AgFAboVVb3A98C+kBjVIphT9I5rO2VvyakzP8PCXa4Rlz9ic98gHAPe40RdPf+8fcqGvc
Y0qLxSy/wUDl4TvFbS7Q2+/jj/7T5URl8aQAEjrmyEOxB6XSXtEv3xvz2/AYHjZuFtc5m42A9nIv
pgEIR4mtP3Bvu2SlTaAsEmhVhbv7LCn3UgIwQ6oE45Xt5CK+EvI9K6TLcxJvTuvcbx2IunnkyjZK
MWuT9bpOaatwwJwnniFe/2sx1AiEdwL3ZKnGocD+O3L0m7Bb+2pO5xUGY2ZkPGnZrCPmMV0QJfBJ
RYNCuTnZBiTe1wt+6NVreHEvQjahzEYIg2RwHDW8CEOB0ULXF1bdNFCwB5bwKhh33s3SBh/rgYmS
fnAfyo7b3hfIVAVATKM/RH/tF5RmkeTJRS68NBbggj/bjI/UuPtPQm3sNY/CylL0I6W5Wwmqlcr5
9n5kEjD+bH1o5cEvP5zDefYWoJ7kWzFx8MY3v4PojQAMQAV62JfoShr0mo5mtnPGYpMTDs7Y5Yk9
6qSc1Tdmr3Wc15viRCvdBLA/CrRA+ErFWMcP77GEOj7KxFM6l+OZUcyZjwB+v49DVfDY4Fg/b3q6
VYcV+2qZDDyLltnIVbzo4r0OxFLohwpEBnocYEK58MKSbGS8jsM+Psa6uPnrrMAB14214oJaLg+2
iongp2HAigBEJXCDsQwZuBlYssOzxm4YUK6OUSYaIMigR3CfNAj4P62PFXQhM7qIt8dPbMeYkYOO
hwSj3AONDwNaObzltxDF0kfE1PSLYw7fBrfzx7KwQsVSwiTBQJCTJiYqtkVinJMCjEXpmV67+BR4
sVFGtcBYqykmHe0I67Fz14ZyoYovByYnIo9zOG4KAkCugPto1FqdTaXAVruFbJLSjLDDd6B1H3L0
/wbO7HOX0gf+j1JuBUBCufaOhIQlmARFn9vB29PCf4eMtOZvIqelHQsRWdcukIbZoKQVJFxVC7xu
tRpO1iUnskH3jjPEzfi6FuLO0OTMQV7I8vJkLQQSoZS4RtdVv+5RclWp9OeUG+tC1RSK+i9E2VWC
nz7GCRzTy9npTX5uF/UMBvAW6gW0U2tBZylFqS/R8PEm110hkB7MgZhYn5fA874ZlXBoXRQ44aSj
gVCiddhZZ5HYvO+3A6+EKNQVGW46dXqEPy/dU6p52lix4mSCQtmbzX5Zzs3m57VxB10vCipeHic7
gDxKRuCWZtrpQIQ4lMilsraR5amU9aB6HC8zmxp1TSZZ0xlZdS5PvyQ7J2jleWwv4hwQEJQyvOdU
1w5lYjmcSGczUbN3WefB/xBLK9DA8xY+xW4O7gSwIqAC1Lf1b1wAj07bCXKbuiScUikUSEdSuysW
fD08mFz3Q8Z2rheAc2CjiYhaACU43hSwG3WMO7PmpFhc2waFUh9CQIUru6mnqUyYRCy1Fj/RMygc
/1wyACO8mAC3DYl7tvCArElSaPQOFDVg7D4lslGhhPoflYLSTSn6AeOTUD0X9enTFrXLNUlA70SH
p4rgHjYStUf/Owj1l7a6gcre4+Ink3ulngzVKKYZFEzz7qiqrCVwlq20ApBc5yDrAFviwgvQ6g0G
NO1MCxfeGwNL0rK4BfeFI05/CPeVmPac6aZfSvaOyhLqc9zyHSItjeG0N9ZYoY1rIgo0uSev/DX2
lj/cLM3TuBwZCE185KeV3LFh/bI4HmHwS9+1u9HtYZMhQNbXIsZ9mZDM+WmxUktcO8498wMrM9lY
6yFFVupSCQeF+NvOqA0dxlv9X4iqaIElHTIMzj2tELy0l9H2bsaW/GLN9wCLkHA3kDpbxiXpcNIy
RGKxYEIlsXEe5PA6Cw1e0VPknRZGAh3NkEDo7uSxFbfRNkxf+jB1BheVl6d1ClOco1Sr9j9BCWys
FsI+vu5N/Z7c587Lbehj9il41RhH2pnw7x9mD8dgNJIQD5X9ZxykXAEfyEKLqU0eHdKpB3q5MR1y
eXSyqBNAhqL/1OglBPb2W+DRc6O8woC322JeI46evds0YDVoZE+Z5nCGty3xZWhbUQFn4rFsBXwd
mRoZj8dHJLCzqpx3tCOb2iOZlnGYGbosaHP8LQvH4shWTXf+NNcTV8Dn4zaqnksUoy/dp+HbOmN5
2B4ChrzsZOdXSzhB20K1oXSqLrW99kKZ4qLhcSBE8aizlhi8xZo26eUyIicz2S7ZTo6RZvYBmPy5
8PFSAcHLzq0Zmrg1TkSMLFbEutsb8OPs298V6RQwE5Mwh4anvGrqxiKZBdv0CZ4yBR1Ry9AChq//
jP7Vm3RW27IqurOsWogvptlSUEHoe1Yl/8I4xSGCiGPW53irn2BORhPJiDARPaqPRNuXtNXtTdLV
w/okFz1Rq6m9IpD31L2ZOADv0oxrnjVHU1GYkUSfIv4R4HbdEXumgMfCJ196QT02dD42iP0EWMol
NhAcwdjOyEPo5tHhqYYhcCpPkHaZd20tgyFmL6D2KHlzKY+7HOrQmxmR90+IIlbvkkc7LMYsIylP
m3EaEnKfmRnZ1QczaLvCyYNEx2C/zUOdt984s73RlsM8D/ohECTIGXSX+4qfajcygJMjnnq/Y79L
bXCoeCuyLEouDqQQ7h5pDwESqQ/XBgvakGWphgt7lZQGzpYB+u/wqhKEH9+aaWid5et9PANaw3pX
nn01HsRG5Xd51Cx1EqJ1SKqFqlRIifhK2uIjoouzd4K6T8iLcF3G+fuPoXlVemKs7I0eiD/EdEUA
tp6Kn84zdMIpgen9tWPWAfqUVDPdQliIRQvOlT4VOLX+N3+d0aKgIJtHvb1TFlp2YrA03u+9F5Qc
8JeTFz8F2iJ1AF+1wxdecAnrSTzoTGCsin4H3Ea+iO3qJ5NM4Kc6zhp17Z1Hc/gA1+Zu0s1wYqCe
hFjxK0OJ9eF6qvBMfLMnoH0aJBQjMHEHhf51NXzud1D9RPqVvoMUPsSW7qIhEYjfpJCfq61bdUp1
A0Zy2ddQZuigkL8H/lcT/aBm2/s+m3b7qR4Q9JAuLQJsia4bvIeOn/9T5wT9SuptCHrPvuaa1ZyA
6Kq4mwhKr4rTWjkBW9ggxIU3DMKYUjMLNiqmyq+D+FgCuqW9pOg/PJJYnmmRYju4djKLf3QNnUPg
Y/ofd7ZVRq0DOSpNZIGbCz0q2TABRve+Tj52XtSwYhepALD4KHCu5v7iUFdWlZQVcS725t29oX/d
rUk+ZmIbkVWfJX9s7LXmGaxewSnpfG9hMus4TWlYYomVHALaDJ8XVA9QKsMksCrn5gMvCQ7FUsZr
pwFlZGOM+aTZyCS2SqieREc6Q4JwaxwpIwmMz5xc+HFxi07pc6e8pxrGf/zATue1Qo9Y9MZJ1HIw
7MRZlxwPyzrpSSwvvEWWOGVUf350HtpfytW6cqovn2uRHf/KU90m1PmtMmPqaEsQDXJLqajm3T8U
5DjL5r3ru6vDDe0teKNF5lt4MGZWStBi5YMk+Qta7wwjN1dQjzsMfJwNrFT/nv7+8gtCpufzbUoI
z+di/Q28vRrx52vnLccTQjVtRJe9+beuYpP4JiLVoneW26u1gYGcyMEKE0ZlzUPKst2/yw6go2CH
uQctrB8C7GPwY5GVXEZt/WV7DLGRVqfvYw+3S1tz1N0/ifXZjx25A/br6nE/siMjRNJ1OAncrxdE
P56/sN82jhksovP3j3TD6pqQyLb2feTg0NcmvGcSCCQPKnxQNzi7PZYB+tq1ohFAl6w1a8PmKeXC
hapCvRBL1liwahVs2IZg/2ngTZmiW+57emmeYfgPjCuafATnVJPgGGgyBKYdZkJuSb3G0eWa0wL9
yDRpL/QSG28JBQ63QizZuuGQhC4JPRaWNqbDF7L7ijm/uQZyN5bBZQnn42DYxtsbQuu+8Qgw13Se
TnzT1i+1ZSz+A6sec2i6qUVTsqpm7nJiCzTK9kH0AV1Tq/TDdpYzEUUbgsOdj8n1Qk7kVW60pWC3
t01EmQeqRYjga7pgZeIOqWiGYvXXoYD/oXHSfZdQElzewYqN92FU05BrmhN/joRWzx4wnmp7PN8b
+4/mC4cAx9ALWvqFYBEmQT5uR7PvPBMNBn8ON0ZJERChFeloTPMfnXBhQu98y3FeuP3RLztBax1d
XaHKOKTJa/qRMrqw8sdkuf1md9E+2CRmR8xHve65g3cz1GHmIriu7MkDS7ZwCOQGzxY9lHygYUub
c+EQf1BtUUG7ayO2QL6YqEycNbYg8txaLBBG6MBwIMv7K/29vX/2RNXsFcKsEKC0Ov2OldrgU2oB
wdIVct8nfRs+ngUIwYR7dgmvqNMOnAtwMmU7mR9guQEpElqhp50LidhR0r/VzRzSYazYYiho0hFV
FZ2fZCVbb2ywgZi6xGl/REO4Bz0Lm6OKzhMvUjur6EQ2R/fsUx8AisLtIHx5lRwM22+NQH5z9Q5L
cmb4044+/k/V42hNH9MBwN/bpEmE/oO/iS4e7osh80XPtJKdF6RrTvOhtxC2egn2ik+Pb0g34Okm
NRVRvg5GrLqgvLiAFrwibC/tV3Lxf6LSRC+wJrOOqGfOp8lOz0rqPpwLy63a9LfRqaD9aTM1w6Mg
0Vyo9eZg7axIQGF1rtA8IaVkWPkIjYKZvCD3JKsXsXyMfpK6fttjdMrq700Ah4t8lH09YN//Bw4e
RbVhHDh9N7Ac4tmhsEhcm36n2u4+0EvCYyAVbJ7Bff/xG94hUjpbzY3we9cZHGvj5V/cKReII+HP
m3mcGMca8SdTIhzPfeVPnbVO4gq2ovBn1N/9S0HRlip+RaDD6e9wIsYqSagHGug8ls7nvA8/Gylt
pJsPpZJhyI6ZSaWwim6ubfEGdXekbkSjUeh5s+oeJW0X9jja0CplA06ofL5qc4D08jJgu4AFZ5CQ
AyazLMocL7dqPL6U0oeV0tvIhB5EaMgL+ldtf089Re4yJ3l9PJ6UNdxpXl+zl56VaZ5hzXvn/UBB
KnJoUmORxb0rzFhYcn93jkpbCsQbivaxFpmLwYEj1ZnuxFymyb/HoEXu/830KAfMaykkf1mFuOAP
pUM/dJBp2QZrokWQZTqFa5Dm2new4zEDTAY7efQd8erDSbcVLkTlTahekDLrb0OCeZz3gtTgmrtv
DWCPfpBRMBSwfrdY+HRNxZDgjluNc5bkOZLlFvoxnFwa4lYhi974vtetqK+cRU9b7z7Z5jXiGf5n
+6eqqhL8sJEj9jvBhW8z2SmWROWXkkHf99airol8OtVeYHRCG8N3q52tyd2tIdFh2uImxJcQ0LOF
Cur+XhzufsCaSetbQZBO8usSqOW84tsWd2TUhaR4LA8Sc5Fd1Ds3bePFiqAx20pTUHtw0nq+dZbB
ZSggug4aFCVoWglb3rzmtyLiU7Z07DdB2UMEIqXyiQ+i7BqFrh9pL38jZKyLyOwtuEuUJh7zaK1B
O31SPpubXJCfPHbs1K0g98ntGu25nZEm1eGQ5mj2qXoOxgGoyXlcS+jCMSnxNVJsHmtfm/LdSmmr
pg8dOOKsujgmsV9Kssjl6k3RMWMrO6s6HBSDahncWrXcvKvLDLpKVQc30EOUFIwxC6cNjh2Yl3Yy
0KU6bwe6EcEayUtin6+VSEGHY4ekOYPNWYweyVfx8BbRIBjmymuicY36WC6Y3EkK9Fgq2rpjvIhv
nb+RBha9ZRcKW2z9+8DegEfn1vMkP/LBwnQfU1mbkCJXNNfGKBqLP60vGVQPswutnvtO2P7V1dnA
Lm1tPC1YGzquxdk9W1970OoLtd+GH0XPH40+uM/PRvQx8hC4Hxqk/sZrFUgYl6z6LWZTIRF1yifZ
yD9YE9q8UfTsRphcmOtWK524CJf/aZaOZf1bdPHubJv5QeDKwb2VDYUgmD08fLmAuy0LCGat3rp9
cRqrmBpiLXs3A85EfiY8H/5ojEKoM29NXdZWJ1d5mhZmIHvsJEsFwug6XWw+UjXau1d0VqiR1SMh
8+ALzorFWfhf9dSKGGhT+vrzVXpo5eK8smNdZ+bF/CQLcEh9995SVEFxesrGL0382/QPb2G9Vw1y
ZizAWTrRvew6BkWAhwFIk44AeMH7YWFxohrg2eU91hYFAU7zdEzGWyV7frzaaqJh2t9HmEFIdV6p
dyzNcfRXI831leKluPO5rHX2bJoy+PHVdsQyF9+j5rYDb210oiYsPm9TqL8M+4/9vlKAnUG7usuZ
J/bum+62bWKEc/JlZSWBqBqLXhSJ4mvasMq0f5BRoOKtydfZVLQuTsloydm1SN5RA1QWz3m1MMTo
cPL6cmchxpHJSfK5vCJ9EB+CNk1K0gNrR0UE5ZqH7WSSXi8PWdsWLwKUBSIYSg+LYCcqJVIcbfcn
sJCxVhLvIqJDexhBR6uBx7I30I6vorT+v2N0skkIU0vScCn095q25/aRcf1jWESBs2CVCtInnGpU
xGbAEYaAdEh7lbcTphsbMfJSpSB3Qcs7Xt7hRI11Qoq4FJtwQMqgxzyM3BgmzZaLrxgls5yxyOGv
a2ZcfYWNjrXHsEfQrhnRTss+uaYAVXYR+xsGA8BxfZCMciEZvzhZTSKzPiqiHWjpuSMjRRFHlLZ7
3T74dibix4WQyzn8byUEwUtlWc8I0LgM55wVF+14DBm+HrfGwWZkjEI53DPZuHy+7vHQ4GQIiiox
7CEsgkjlf92sXocFpNcFL4tP0+UnjhDa7OGHb1y55d7tMpIp++oCbwo3jo1K4LGfSILicm0bdnrF
y8/dd6Slpa/jzExqwvHTiPUt29E1YPuxGJ61HWxNeFOcCHXos3fXxdX54eOaD7XwPgSOjksajJBP
Fz7G6DicWlxOAa2tKjJOSjFSMWIYt4Hp1W7wdwD9QzW2eC5oSaifhR6M9+tFfHKdLG3tbFsGMSwo
tLbAJCpBIRde2Sog+3xgexlwDAcCIAdsNNJPWvZyHc/7bpeXR41zZh62ZUnYyQFSanaTNghW+F6q
DADFKNma9P+I3wew9evPW+sLrQrdZEbuwfFRNFLvgrMKQqPiSE/nZYZUYaIditsABu2mxszbaG2Z
L5q/k0Cmk9a1HAqbOI+V3PPAWa7Nbg3OThOA973WrVjn/QTm99nNY68mQ46p9Jf3OmUtbNw2EGeM
wYElu4/fpfDRLtbml+wEEu2aa2Vls6B0B7c2BP4T1aZh99Lh+ap4NXK+6eLkQY1cBup5bUQ8J9ot
NPhMHtRqMWBdbkJlyYeW1BmW6eA0hZ6jJQ5rf44Oj0gzBJs38eRLviCW/0Jn3a+7tMKnp98zZg9y
rLSkUdsF92SdBcfeACRgCEG9Nq0FL3xPXG7vbb8bId+9/RAEkRuve8L9jKrD70m+IRE3jW0qbEd9
uiTCVDp+55tKVk0YA/tsEFTT9/p64Ds5Spmur5BwwT7InQEWD6onkmjgnE2us00CQQcp+M7E6mzG
ZKE8+hpK2CQpfO80Z92Jd5lbE/LFDqcuD2NSfw4eEKlJwHa5Dom3T+Xs4p7XrgbPf0i4sI21Y1pS
feq0JrxsUcgoTNykpvaF5ha1QaJqMaP3wjYvuFi+FNHzeR3UIi0q1CJCkE2akP0DcyJMvPLKRQGB
p8TcH8a7ZnCgVug8U3OD+xeWMnTGs8Ubu6pk9uwt/tPV5solmMs+EEUiQRtJmdp6qmEpxaKfShHO
j77wx/mcf19DPGCtkzMadpNoez0zf2BGmmDcRaKG6x4b1hpQXRHfGLJUjjfDER2wPVZiF6LepDJ+
EwMlmYGm1kvKDVKC/Oi61FUr5ss2sGMZMfAPm6f+Ier6Xi7NKTxFrfklimIYcl7Zkxihrj5RZGDQ
5g4sMQ88/P6xzXd6MbVB31du8zY8WiaDi6M4BNYWJLNOFeN7fR+eK2CnSXprWXnbuCl8gNjQhzxw
ZY39dSzb4kmf0FlQS7DrZ+UoY/WhoG5PrkuYwk4x3N+Hsxj7kMBgVhgKLtymRI9ZrOIsh67A9kc/
dr9LmfmI9T8nLyAXTbl9CtVHd9La6La4wEsfq5KAXKYx7ZHlskVcVudIu+ANhFzDn6NZ0+GORgWi
iQS/Bs7I8mjU/8g9sudZT/1PLIR0q41p3GOllWb9TbZ8kJgk8ULGJXl2B07bZ6cbigWHam4NjrSd
CTS6+AaQGd1q2D2KTQ5xVTAMEqziWU3Bfk8OTw+V1UeEzkmZV6eGzrb73xjwL+9WtYDw8B5cquPI
Sa20K7BGAWzqY7opftFGPQjs94OvSzibLjrXmpkImp1wflgWYDJ6+ApbJmS5efplVZr9asmjtCDr
vlu9gE5luYz2lkcUFdHIRrNUZ1OxJ8jVoVQMJDK1woLUwIpP7Ti7HD76ju7S+5eEKYRqTZWDE2c8
A8MneDpCNsGE+Fnm2QivTOz+3SiLCzIyZ7d8ibIrdBCJJc5estefto6CkMvBDvbUOjyDCLS8KVXs
WO4Iiaom723SZjUN1/Z/zZiGSR3kPU2xN0wwJh6j0lO8hOk2YSu+1cw702wPzQALMfoupc5h1zC8
L13/X25DX24bva9D8/0GGWRo2soGD3hMfiM29CyNbvhJjeqHC7WLXhSWnX64kZUK6a0aFl8i/ppg
VyhJ1BaNW6Gbm08xMiN/oFuQD8mTW8WwD57NIWrljChs8zcBiIR/mH3kRpgH6yjbhsdLJpAtxs35
eUuDYC9Q7w5bwfs9iDtxLaaB8qbTQs3MwXrkooBofdAUAAwAiyEtjJk6Rar64BUFklSkIRNZ34J3
oKtKmLZ0ZQSY09wag1x8pTiZUlJxIR+2zZ+h2n77U+x9hKeaAJtNg7zohhSt7YEOl3M9BGiuVuWf
/39lvdKtPIbLIQCc9+oRJ68nvnDl2qR6zCaaGWtv1B7FHzUs9YFWZeJFNw3A7mGo7cAa6CB4xy5W
KLPyXdM/D5FCvM7SvhvLnAMUuRqtjZnaGJbzHElj08JO+xg7hTtTxPlWjjf8lJDZB+fcalOqweCm
+boSRlyQxTKwKlC2LkOxI0Y9gxXBc3WC2DZ2bJABUo9boI1zqxaA9JnzJxbFV3iI/2ZWgWx9ZBY4
rjxEtlsVhMnJvwsH6gxgMOihgbMDaZbnMMhARRueSSPZ1aLa8tDz6kHZTJwIqjBuZ+QG4BwH+64j
fkerD2KzrBQm0MSJ32EeLbGS5SqJxNrtTmbPD7/UqRNmDbcmjDLy5fFSMIwMR6j/AcSbRDz174bl
0gXqm3iRPcHiMCM3Q3qw5ScEwLpRp+hPt0uusmsw3F6NuKFwbd/g1wmet9JRnOy6pReWQ2Mi3ac9
XhsKwRiEQaEcXrbWTWE9oH/Z5b/3vzZRRgCJE2cQfOyRLDrPyh+Pthz1WzAc3eE5jRnScjJpuBw/
M5h39OhRx73pJ80TYeTxwx0nrsV2ITCMmJmIXBCN+3+rdwvYEgVRhYoyOo5S9FVi4yUgfZhBn7lU
WIF6haqZCN+4BrOMOcvkD4z+0hQbFl8Hz1grLTF9J+RaA7qRKhFOLqw6tX7dupFaf77qWw1kjp9R
oJdk7LTviIGO2JIS9BEIDN66tkPst4cVQdEzGRTJ1UBIemcqh+G8imgj7zXy572Ga6jzkYuzp6Za
J1TRtKsmaYTHLnZatMp5tAi/B/bT3RiDZ15N+GR6NJq7R+6b1FKYVB0/i2W007z7ZJZGhKiZ7lwv
UrQB6DMn1mUnh6U1LMAYE24KZp3YGiiqI9+4hIaquE2gxabyB4WgLKxEfzhJKTdCZdIN2k6FgTAf
pcMxsDDoxAkZya85mEtDpFwx4w/htbXg1IxzluGyy1MYuFLZtfVrXOESGz4AErWSc5wtKkL9vDQz
t+Tcnxb1bMoeAEzXAxo1FLCWo+wF0dL70YxEWXyyKhuj1aj//4eojQebxhNGtK9xOLs+FBS1D2J+
hBQTmOy19rCODRwWN3sd4aM/Uo281HhITX4pTSoE/nlonwjiQF1OfZJxJ+Zjp42KVV+Uy7/NUJ2v
l2ujNb7NTzSjYl7O9+aybermNBy9i/01dvbge3o3xUdpGpYUi/17dj8xyIbDuoiYCY/yGaLUzj3g
rrPNXLiXgypTJha3cWg46hPLHVzO/AWQHo35CPWKkVahBJfh9UOEKnFi7NSgBIiOpyTskJLIJzpm
FX2LqBawEP1hOgZe/IEEvpGydeMkm7moz3NKsL8we/nuQf8GUkfi093soFOQCujiCPCo5KqFAMTe
PqQRvU1U3ikaputHSJF/ouR+45wkqg9lMT0TZ0Cs8O1MqKopi6NabQfLPiQQHBix/bUzI34MM3Dp
ZieoY3nM4EPECngbnS5tgyDVK0yLE8vQDWRh71ek9ChI7u5g/R69gjgcN46B/V3cnkZh5Drioe1c
VKmYAeSm4lRXJUT5i+AgVMFBOxkQAHEoPBjxB52dwqBJoy2Ip8a7PHnoOItJJVaLdGAy+2VByhWW
vsODrP+88FdXNqMrjn3pes5+95jF9c+dFh5w1+rHgyk8C7w2uS5ZZXuZqeBdSSP/se6GDsjbVTT3
0ZNLU68VSQVVzuoxIy+X7gUbDW8kcYwii+xG8fUeLzSKDC6DQyJwC9L6Y8NcbAiGmnoxHazl5mHJ
4v0DgOUMKb4dk8tLvlv7KpxX3f6R8squIJjZmdM6JI4Zw9T9L3scMSLSMmRp76NRfdgIzdY3ThKC
HWlHKUSCsMbi+RKqZGmdsgmI1Eoj6JGr7Hv9jdAOE+jNY9TtTPfR8kX0sqyGtf9URSPcBdZjkKH4
FNNm5uUO8sq4VZa6HorJQNTFqGUrDlCcA4+N8YvUoxmr22Xf5Ph6Kf20bpT1gxu8WunwNEZ3SeMY
XUuqf+xWsFUm/f+BL3Ihr6bSFyoXA8Cgva4QhUw1IqmyXbZvIsLkbveJKAh9U1KuK4uUFK0HRKVJ
UbTOQeW6Pryi9nU1tw4iL56q8N0zwMaHx4HjHIQ7u3NSW/yZdif4Mivee5F01t6ECSTj1OJNPY5T
iwGLBQeonJ1Z5EGfZnl6tfxwovF5JMsN2/j/kRfg6kijW+pIIhaL9w1x7ScEqdM8XUnk1rkz262D
I0eeSTyvjbSedQkeGbU3QnWPnksV6eXSztZpxeICR4ajAZJeDltaE4Zu0BLBUiahro2eyqR/YpoT
BItBSLL40AzE6bIvR73cyl9wdQgy/9oNZl1nKiz2Xd9dDxWpK0omzxO6m3hEEWiaKw2ypCGIM0yd
tMJWEDuB3f7Kit3Ps5WdpgSluhfvtIZ9F3PKZevb47kc7UiuEhGOeM5innPxgDPFbt7SeWGvhoYQ
9/tidm3/1JFFqfHtwVuiUyAOZyb6/AIRev/fyC0HOoKoqcZoxcNVthsVnJ88H+5HAar8DJwME8QR
VaE0iUbvQkBsKGZAd0cwu2KtMfw7/rwx2zNNpAa3rJI3/867WaqIO67EK1TgqR7AcpFVCxbwmgf8
1m+3EAHZQ8WKrFlA8aQgEuPWRLgh599Q/iBjvb5gM62sWObZGpQ76Cz1V6hYLCszytDuoIySbsoF
ugv/zS/As6LMG/fw6UYDeIqQrZFe/jHnT9ZMNFlXhkQpmGzOhgcz4PXGk9qp0NOscsZKLMEmruzH
pfWGg1NN2Tef1aWnXFpSBPJltUh9P8j8ZSCM2lymrmptE/wzxrHSbXH1XW89g9VBTxfjcWrUs/S/
/0PAX0UFcHWIPqdm4UJY380RWdNWH8h2LqBFtALiEtyobpe41nCWSuR4XkPg3k+kO0h3LM5sU5LW
kRiTXiHe9EVX8Rn9VI6M4U87D8R3PukCYhxY1uGX8A90UfyJKOZ7n7kL26QU5UoegZHau4RMFswu
dYdCamkGJhrGd9+CBTLVm3qURXRzS9VazidWketO9UAtuwhTsIG/ZNXzta3RQnCM29KCMQOPnMqh
zw+W5suPQN/GR5FSJvj2r/PUsthgRpL4vQOXwfBGqdttRch3QdEdfHXvkmFUfLZhsH+zP81CFWUF
w8kstWzUEXbIxwJMhHP+mxC3V/i7J7CkOvudLGYxXTSkB13w65ooYu6HE+7dYG9jE9VUx0JWUknj
w1bfw7kXY6HYS/Vb0zEOD6jggcXsTSOiazBHFBpLwOSg8vzptX3eCzEgZb+GSL82mHqx4xAywVD+
75hDQ3lOnYPciRSMY9BZhH9Yz3CAKva3Vf1hdzu0uuXcTLHWBykJCVx53WcT4SAukTAk0kSRE51G
VC6C/gbQqox/vq7qy3l3VkJdRDeodDNIIk0jCLEOeEW92DxkBiC0BYGuJSFx9lPzFGx8D6eVZE5v
8vPcJ7UoTLsJ76PqhICX4btEF84f0n9JRFa6fMeWWM328hYUG7Ol2sus172sXo3EFsq19NCrS1L9
jqFcBTHjfATHDw1p7G0AZHF2X6/NtE4cD4GKN0ANbaXa04dhcgqpeDosU4ptM0xiOUvkqKZQTGcv
6M9miNZbf82i0S+gfGxzP8mFYkmyZkc6ThuLoyRjbFrdw6xyrM46GmfSbQUHT6Kn/XjOiG6EY8i5
IFWVUZChKePCLmo1iTQhvtLCwRQzh3p9nfllA8fWMqlROCV1qeapE/wpoDrcU+9a9EIdaAXS5R/Y
JU/Ly+sX1aAyAkYzgDgCvC+75hScNYHtsxTaNf8CWeexQ+YKYyfpdq+cRIjK376yQxlXZ60fbxqg
WexG3cLyfs8Du2X4YEeLlF/naVZQ9caYPHua2TNL1HO8v6LzgWmFK2ZOgI2vnp3aTnuEVx/ln0X8
JZrFPK6UzmLPF1lNlxWyILpRj7/CTxj4FhdpzQqKTj8IJJdDY8CHbxKWDKZwY7Sv2z3fun6NQV/L
6ogzU2WDy0xlpgQZL8bKOTKldQwH05rhx8bfEMIGHLXMwOZmpzBDsMPA6OtRag+r336IA/LWn0FD
9qJ8BxzXDUUuslc/lJ5uPhWy8Ea9LEj6FW+jDogkmvP9fgUVJJElaFiFvWJ08v0IgEkib64zj087
D755q/4fg3AinVSgr+UmRrT6Sflh1afAZKAxotJDCUjcNRrpTcmFor+BH8aEE9uV2Al1v8Ug695b
XsrHsTuTOC9wmsLwgxRGu/YhrgcbbDl/wTjnJ+0ejX3LkM9rU5ICjQW0vw/ViT48UEKuC3kf07Y+
zsR5/6sJV68qWFIZf/mmzySQINN5a6f8PFxsdG83aPQOTEFMAHFRrmbhoh/aGNmraz7Sb7FcfZqj
SZF/+kJeQ63DvP56ueRgXHa0qlbmQjtgAmd7LY8dq8fY9tvMwUap2v7O4VORm2his5YJ4P+44TQk
2MVS8ivhN1pdjdLEDHqOcBtbF6ZDdjCg5XemsWS6JtFljW3qxmedjNzm1W+PGQY+ypkIWfdcKACK
V7hHHYyU94tzjMh4iv8ra3+j1Txhe/ZwZjOLeniEF+FMVFSpujZLT7aKQNZ75IDMjyxYSbOtXh/w
CYqQpzWgqScWmYUMUBwhEU4Wqis9ySAmRpDGK0TCbBPTyDQa/NgXdum7iA2EH2hCORC2u0Kt3k/a
BSRR9RGgv8LS01hk+OeW1/EF/HgWIIWvxAtQUJJ7m3rSonIvRsEBXDCXpUicq9cI5SS5/KH7t0xA
A9L21oPwGg/3ozXog/4JBURO3Vzp7XUobByLuK5rncSAB3p2oCpsSPAM7VqOvf8LQimu9Rov/40r
wXsd6Yt1qUmJ8UbraMwMqJVTiyCvsxXkDlMwK33/8525x80NJqSZM+akyGngVeITejy4hweDg7Vg
MfWmxAgoUaFEQQ8sMU+YIzMO6RnNvofkrpn8OTtDtKRZ5wY19xPWhD7111r7VjsGpXMp4uIbkt2W
CQh9fk+Rga48eAtGWHRbfX1wHsTPbob99v4fEUFOIS3a5rmiNoq8sRmow4L9RgOoPXG+vqiTM1Dw
Y7m/vQ8PoCWVvu7P/7fqEiGzspxRygLWHLxgZUADsS6vTf0jWeEhWqulojfdpTIvKTc66IROey3b
8XiUQGXyDJbf66dD9eq8cRevDBAk3DLvC1F95QWktav1mWzsehIHINMNk9g4qWsVtrUAQah7iOPU
3t9JzkXIdFmh+zKEmaA4CWDSo+LZQyehn9cAOu5KsYfB1HWjfN7BuuE524SVtHDHDpZElnDB/+/U
rdGut+G5tHF00m0EX+WOpHq7os0waJP9Cv9VfrLzNE5qQx8nhCOgkqNQkAheIOznO+C5U5WS+1a+
Q8Zac3r57o3cnc74jATgWsK8JsF0kGz0B0CvqqhACsu16bykj1Bo94aCfJR+BKCEu0kCfp+W2T0x
/WhSv08QX/0wIzFzRfaeEdIA/TDAub3U44uUCMqZtWJDDZ8MFUEWYvMfVWbc9wmZRZzW1eDfrAoO
rVcouQe4hFPnR6NyOYbVCTmYFemjYu/MWJYDVuNEfkwbO5bION1AEYEQDOXlHWc7A77Dk6OYnjFI
D/Xoxs1UCprbu2PaSlCy1kIEf6+niQP4fwglDUvV3e5CaLjzxxE7yG5E8aa9EUSMPDGQTL7t7FfS
1rULsoloYhLoCy+IrHDfXiqZFZcAuWTntR8HD4qDlhLLjRqcsJ7z5ZycAK8NM3Uz/mUh7ybg3XaA
m6vlsjXZDZ2xdeGnK30Xtd5626PvTfCUZEySpzO9DC7vt9So8liQJ7zRHcvqaT213tdJRs5xWYMZ
qg8y3VEKYnINpjbk+lMRWIpK6hE6lSQXr+/5zUoS5H89YJU8xGMdzTJOvgyLHsz4+lkf8RgBDS/n
MjCGb80I3G/GtyZkij3HecQDtBOuxG1m279NDx8kBLUj5EAMY38Bpak3LWuIdv7V5Kogokcmj2cs
Pu1lXWlXcdxb6ry4RRVstIla3YzNs0mw5tz5pmqZewSWc9FyXVfmSUt76vtDXGW6x+pSIzBO6mwL
mfNVq+dvKs7XWfflVRz8SfeUdrKKlrisoefRH7VCMI2Sa45LNKT9djfOvizhwilDlcGQJcwYii0w
Ny9IkULO9Rvoe8hOl8Bie6qD7W71dJpxVxw1r1ymkaN2Yy7v7C297UWwQFj/B5Ro7FNU1KMN65kO
4+L3sCeCYdqLBOpE7E/Lwc+myszTydOqzkxfaFWxsIOuooDNypnn9TJL4/sN022lvALj2e9vvjM3
e7adfylOxbA+l1uFgYn5o8Z8ZNHmtfmxkmB6K2+2Le2VnYPJ3vQFLld4B/kaCER9FkkrSJWO1hsq
Z94CxjTLm63Ew/+kgyEfnLtKn3y/Wj53dOvoRInvVGcBnIIPY8I8CpDkgu1PrxCguUU/6fdPmz4R
vUvA9+Ypm0YVJiSY7IEn0sNZ6z+hzKxKuj57xZdySFcN1szobaIdlMJtkcPT/0nwtzjwH3RO/Bly
R2HJFcOeq5v0FAX5Wdwh6J8LesJ5oUXWjW6XOUPlLVtuTmDnCp9sPdvJBl1nxr0XeiDqHPBBVcKW
UnArZLaAyM34c+XRb4uodaXZExRhfo6dS+ds+w4lcSmBqtrS5mjd0qsd0eglsi4XZEGhwTU9dGCy
RPmkdAellLg8p1MP6msyoUgRBRD380gre+42+pxkoqX7ImBJKRmGMjNofPbpvu9rO1cMuWZP57UZ
HQ3iJcJ3c+cxAzH6qATsg+4H/bkU9+Ac8+bA/kPn8Sztrw9fIkofCNWFPoVDveX8Ur0KPoaT8zaA
IqNCQ29ln4WLJtODRUDskRVcvx+2Il1VnyvaLWOqDME/wNTnrllnaI+bjw5zjIFISdlFKuk40LQN
i+XUMvjRvpIi+7uCeVui6doxy/RcGXA7GQH6Nm2vOj8wrvYPYKHIm501E3C6CCCNRKj5iXi7ItSi
mI/3tBLeluFOKWMhxjVvlrYKLaiDteishIyC9dxAuJ7XXjcoC5rUmya/fSmGPog4AnU+jAIo75Eq
3NY6ERNUCVRVRrlLShAeOO3hynUk9Rlybi7uGoA8YicZ+t2Wjs6WYFRubYzIZ+TVVlv+PUyxlJZK
2cNpR3DJiPK8gghbNTOgcvimVRLk3X0bPOkjGCnYqTKGJ6/exEGYYDRDtA8KBcadBYNFW4mB4X3z
eMipP9qEacaF3e2rcvEfu3cz5kUH2Oc7Kny8OaOBPQ9RBYkaeF1dI3aNJdG4AvdwsG6pM495YFW1
xqQpNGz0MsXDCg2Z6WJUdUK5saZJ0LLpftOryk/q7fzqeIeW41xRTsj2EofycEtUFic4IvtJ+0S2
GZsbFnichAXvAG5kExT0vkbu/fOCgiyqqnJ7SBUiy8URM10PLX1/CIKZ+m9xk5QaMxoYPi0fI7Cy
Wzt0kg5/tLNUDztgOpL0xEs3RPKayodGqpzc2pF1zMiFBqv3aOAFMJUTMRX0YZZezui1FKm407nE
Mx9qNzg2mFSce3KiE0lusoBgPE4A2nB/RB3PPBO4xjO/E1zmP1bpjyh/p2d6p8Zkb6kFixCvJjnr
NTA6ulFqHK8jOWIwikutbGKLHvsVCab/9m3TV08qy1rgRvXK6wAW7zwOZcs6AU6xPYpMvx2ZUyZJ
0E3saU9+Yibg1ftj/+SyiUrGyohVFPyUXtEgNYBgMmv3BlcjgC3TguK71FPcTmc8rchi5bydnCdE
sFpRz6b3kIjOt0LRHdag6q9tEEb1rkpzW8bHmi5VuyQZGrW0L1pEyrWg9wcHJ1jRT+Iztgz3gOLc
YFlg+5DkiaNKrZweeGAHCiLcr3Wf92Tc1hqR1Vz13JRyamxPZ5N/6/6eZcQ2lvGIMDhi/vNuC8yY
liFu2U7QeWwAqoaPHFPvVorBvv/0CcoGEANjT1624xLm8G+6aDa9DNVPcceJ8eh8wQZxB1a2sjpf
b1pmhRYnwe/FvpNy5SEWqbbUnN2ahNTANpRG6wPJKf3qhAH/B6F9S/fMfeR5pSiOgLrl7WtQE9Mu
pg6V5yfWWrN/8hNRVmZuwFnE8Ssh9pJ2CZBhXA1PIV17UFEUvpe4V6YxcOhs4GrxEkBwXGocRavz
74Ot13CKBZ/JJB3W6mJfbtUETcJn53n8jy6ymrBZA8KXVrk/LHILMC3WmsH2Vmygm8YMZKnlrETN
w/QREYDPLq/j5zy8UTV6k9YT9/yOjcHwZg0HbNaamTN2o+AeAPyXY7FpbGqH8tTkIXRkxIHpwm/c
NSXo2okKAqEAFV697w6FJP4cZtiDvXSHf3TBra/idZXRakjauiIEyQa68Ov8kUloby9uqmKahY4M
1vYm8zfq6FJkep7ZO2y3/1H8KOHWoMs8MrsuT9IPiJLpbPuZpHG24iTOTUK9eNmMy4Rkpzd6P4ie
j/DHrG3QucbZo0uqTexjAnS5stMfC71T0Tft7DIlOk0ojR0UnJ6bQndBCon/aRmShPxLZ9MxZGku
Z5afg87cVP0blfGNPOUxH+ZIrOFtyivC3snTKiojI06wKvJB5EF+tp6dQi617xADfTL1KmI7l5Z3
0F0DzmkkCe2ey9HhoHqJr+tEKvs5aMlFObrQdkZuKKJ4cBKye1MGw4tnghZw1SpdIHXdLG+6fxpW
79U8CHuGjfAVA3KAMSmJVlti+3eZGtPmb9QCi1w36G1rrRfLeDb9ke7NeSYZTOdHX875eLdmVb9T
8TXK9Njxhw9VLBeEL8b5i+mm3NUuHwB0XoiXKcJYxs7iridSiyue83Soh5QlIq28nDHbfrYqIIa8
jPnsY997qeYw0e/Hmh9m5qESg9CCJp7gpRq52/YljNpot8pe7L7VbPiKY3w6e/a0g86iUPpaBgOC
sJvh0coNXcvf9/MvmlbO7iLKL2i5HoYCFP/pX7so3ublQZF5LJP7MzKudnbIg9sxYp1WNI9DSvoH
UPLZG1wkBFUUSkRRlvb/2gcrJnAFSfiVCKFvaR9Gj8ZG+TccyrCRcMlvk33FRsL3iRU6TjOFG86w
qHLwYSmLbofgWD4X+oN6JqaGbmbRsS1FfxA+EYQCGQHZiLl5G1TPEQTDmoYnhZ8g8xGP5Hxm58f4
7qPxymM6Geq+FWovf6E2wiELuPC51nzLoq9Gnx7KGdX/MAKiGusX9apEE45ZMLr/7a+eZ7ToQfRN
xqh2PZu4uNsskeeG4VB25MFCyyrBFtUCsdNqSeCNZ7eBP8a49mzopT5+Fs/YCANCB75Ldpqw03Qy
FjqWE7bQ68ZEDmu0XsltdzKrnGs7eajuX2hpwT871bUhL/PKvPPpfSLNBvhMTAVULkK6Tfh9SU1S
aB0wvaBY8p6RFy/x4HPFqVQJYQh7IlTOySa6Iis61L+rPw8hk3jjy4wKfpwS26z5RCvS6DPO/EM1
O4PhTPz2PiClM+wWutYIpYxSFCHW+MoRUl3pRAoQ10vJziIxg8VN23fagrlk4gG3U5ZqB/M9Rwoi
p9K2RIxZMLoYLyUv2A394j9aPzqMxUV2kAgYOZRpNFIlyNOFou1FHjQMK90s/II2XSxAt37a0HHO
tourCWTrIyHYFocegb2rkJQa3zaLT+tKCIcXo3qrxohGWAHv+O47cEZ6AwohqipqAwTjszcioZiD
mxYMdw8l+hYsD6M7KLgddaXKXauTc7xy87mAuvRMe1YcYmKBUyn4CK49/42i3dNmI5qf9VAXiqNO
058lghTnDxNWpiOt0Zr3u0xI53/aCneB7tVG71esZ9Oc/tGfE5vucHP17n7DpdbzsbSU037XyIyV
vMsA5GZHmUD0vQxMD5lqtDBZvgBoXtsmcRNYq7jzWYnKcC8uY77QOy53TKwK6RZqBxwY2VSVYoqX
yrUpOOkClR8NSwVHgkYt4ADXaMq8Qb3f1kCHZNZ2clBVyZkdlo3IQbLUvOZJQM8pyyD58WMrWU8e
HyJ2aZM1O3cSIs4ybtZmGDGdLw+3LT6EwODt2nB4DX1G0Z/70bdnCQyCaWQM93RF5UwxErhtu2ss
WWET1+8zCxZgTagP2C+d+JzS4e1SV6JMtWB3D4mUS9pT3D4nGDHl9Y4CWojS3E8NiqHB8p6bya5D
ymc3PxAEa7y7yTupTHz6MijmbL1lnT80p1lkjcDcMItcs3S32XQMrBY9hBr0YdTcFqtzDrr4u5NU
FMjbBN428M8DdskTNRqzVyxo9UxJKNmBZdMbd8nD4P95bCuQF1KqTbQYex3RAY0jv+LXqV7On71w
wMLLcTxTjBvYXln8drJXQ06rpC9w9+KAr3heyhzjLsNSYxzL1MItVyJRxDM16RyjU+7uNZTEvGo/
XBWTKd93WnasdqpaBP8KErbSWEDr8w8H9UJMV8In6eGR+BGc6WktBIU2v4/oCS/L57cjBK2npInU
8QcKO1zzHVQ67LCmpn7zVDwX3nqsZl1SJGJ+czbKslA3TA3Y37lolGxpbUi57bMMbC2LJ/ptVvf/
t9D7tv5dpzJM6vhM75TkRj4APNhKmTthu9bnemTBNL+YDpZFGADQFr8oliftFiiwIXhSBbSKgRLw
jl5c5yuts4qkUVaeZsMlk9CbUml7fzI1kNr514sgF/OtIibV1p3X+VwUWlcB7E9W/w2Ag90jdVRK
8qX2UZ88FPU34gHttf6TdO2EeC04+YTFkepctvmM9nPHhKnRjUMMwCUC4C28/YGACEWHPPKZa0aU
P+sNzndWJwhNitj8MPCMr1cFlHazkjmQga+i7sxern6VFVaAQOoINwY+RDzQo/jFSt88i1TviYkL
8G00orbtd7o5VrxhPwKroaNlHdsaPDvJznp/P5rGj+pfhhsQiCNAo/V0mCJzs3vZiMlNW1fckTGE
nzKOvvfDeNMespA7YF8hsUuSs54sY0uSJByPnV/RtKZ3LMiCPx2dpK007AHpX6p3v9Xv3WxkMnW5
8I3PPzeRyatNvRciXLYy1FDSs8jueAr6l3Dlzfl/0z3wNMv6aMvbiG/gFLN6tK0cTWtxJOkx0GDB
iqp6W5jzir8ZdJjsPWli3KxK/PkubxGZ3h1XpzY0mVFIYTrQSO5VAIi5HPohnXPxzyVh7rX0mGog
GYv8TnL5eskMYdVxT6W+8iZ2LX/oUszJ/fRvh0j0QntZrAmSP2fpd0B7849Q8tZegG6jpa6xNS22
t8nS0jzveVRpSYnlpWJWEtt84JNMquA0CUP58rp4gtc4B1JloNqK6qwzGKsFMu3UJdXNyZb2wZkw
m5ddoForH7KhRN8dC5A4ZyhmWlCs311F4aFo6AHss5ysVa3c+fZACJzlFzMMag4TCeFOFowQcdNR
a1steIZzVsHEwxrwsqkZCi+UPMy1kcFUcoqyGr4xs/0zdPhWd0s9K8jartKsxJY4wTbcCFF2Fn6l
qyFeQ8Bj8ulcQ2cdAj0u28szUqeRfoFeawEw/zxtt2FV0guBgbt9uxmYQfP8WeoJnrTwIFfrTQxC
wBj9Qq15DlZsuUkocYHC6Ka34hozarRrzMETubB0xJGk3rOHjpawYbXtq5gjwqM1PzH7HgiAdfL+
yP5SrZCEs84H2ecY1FLApMtKW1Wee00v5LSmxgzIKZkbJgGoAoFbdYSq+z1kcxpNpZ5IY+GMa5zr
ygkmZyPBbPBJgPeKVXVBZQqyNnmjRcap8LDRDSo2v8fMhiKUIeznXaOAXDIj2+3PXf2+EViySCEp
/Tx6r7Z6x6Kg0c65PINaEuwsRwiKu1hvX0SkKWf3zTLq1AzwNX1nS+tW0QUAAv6A3lTRBnYWlAqQ
Nemujle/kxN81tSbKzAQm+V2AEH73Q9g7zUCX7kh4k713+HKxN8j+/Dioeii4SHc81dWLuZHoc+k
AzP9on3MXXxrNbX2S1c2B+ZiMRs7OlJS5iwvzwSoHiiLVjJ+hkC3k97FM645lX4hOmIAhZhG7M7N
YmKonUDUz1/ZbZ8IyWEHKMOxckhB5o8R3kALgOGuxEQOe1Yzr1Am6lEbAVVs/DYpA2TJKGdTL0ew
PHdJnM8vh3dn2KV+wyJm493us/sgFYEyifWEris6OwFt+f7q8jTN9M8nHUwKth61kW73q0kLQzuJ
TBF4iVkcmpbk5QixGqGeyvhFkJ6wBa4T9IwECm9jxUsxWa2jHo7fwzON3kuUVSxsclBmknkfBErr
Ympc8cGzc+G1dg6nF8qhQSSEoMC3uLB1ifIt26WC3YEBn7vHiTY4l/ypXJtMk8yyw8UQO6GPOElJ
ySdq3UdPJ5cUQnXBXzESoWc/JCkYpwjyIj1xayv7W3rWkYzvQ+GW/CG7F0SKz8rd2gJm8g6oHE6Q
WwuVqK3gWunXMbEYx+84Lu7J+NYRj1Gjs/x1750pNXgO7BU0on98fGpQ5uGvzIU+9QZwWgZrFywj
lYzfvvbCSEDrBtMmXsJZS813cpFZzVVJ9w1qpYRTpR5ZvEDGL/S4gRfxJ2P12YgfAc9Bn3Tba82r
6XTTRhIWkLUyVa9Xd1gcw29qWHXNloDJIaJiuVASMhr4LpmXYnz4jt6L2rMmVurqAEhafsqCp2bx
bniDY/oIHh8BFFmx/wWY2QWcLj//4B52XJO4a1t+ICHDCToEVWNc+TKbIYBO2J5rypXjNqPH/vOj
G2LKsWI1ipVG0YbRe9BTvjqixCSxwFoi1Bgbmc+qg28HaWOmWqtR0mpA3QnhfYwRz4yatS8cl4hQ
nDTpYCie/wwNcCSYpqM2FekPt8MKHGh4G5ieN7NmLiCk22Kl66fhxsbL6iOJQPXJBqsMoFoIH51D
wc9Zpy/GosyH3vp5l9wCKIcO+n1Vf22G+idSuVde+3ha+bXykNSdagt2PjKXak25lnGlqP+ARqht
ZLDI8zNDcDOqfabxAiY9Q3712mHFCZnSjVEuE2kTGBCzbo9gjXbPAqWxO8hbTuZ1N4BigLy5biuc
vvtcsc8X5Xey4zJgrI1o20i7hWOtC9JKESXBCrWn40m9PL7hU3kFMn7gXF6dBE7tW7abfMkOzQBI
I8vw3m2qOui/q1SPk51JGYHVAEuPTF8Bf+OxoqDaYnINn2ylM155M4NEVXeWiYORg9oJbu3nbL3U
E/i8UeXDpAGHi2V7R5B8scmPbCJ02hRuCYA810iac/xtZhzEA0N47YOsgCq6VDEY4nHzYVTRThZa
BBcOuzacl2hpOL1Cbji1GUMXJNlM76H1iXFX5zqUe18FAyKNMNHu9OrD0jHRB9mRW1v94EnL2KRl
wvycdPi5n/RvXVH/6jHwVnFmdBqdaA0IF5DH4eC9AEkLTpA8b1BwFqeV14qPHhtjYGmAHzg3I88a
xgKFD/Ho7ITJ/HscpoVyaRPK4vZaB1cE9RKsXI489bwW3RCtxLvuOl6/u9ZoN61GzJLuVdAWqP3T
p/k57yUKxti1cvIu5N26FuRp+szKe7PtfqYZ+8vJDUK8sob4puDvYk22WnQ7tHB2lC3w4XgLg0xh
Bifr8+CQQKe9rgei+X81O4it1qN9EC8+w7zL03cxXZAkP/2hboyzNKD/GT9yxDBBvTRpgFfUUYUc
INE/JoYNTtb3K8bEuJT0DIMG9OpRgetojQydY+nL61NpWZwFeGgSi+GcmpDBbX0KZC8XB/XgX7vx
0sjzPbBqqQ7z6gRczNyA/ZbBle4Iu9tI20ou+TcxwfMcuZ+8KtHF6rWe+J2WWn/gHFelnOXoRadH
nqYpUH1lIXzgIXMRyVwr4tVM7hNcfmZ/aI/3pJnZU7z8zn+xeDsn1uJ4kW9jAQEpDUYK6eH0aKM8
G1EpCPmsLhs38JNN9rUBQfHhbYq921qosPPyHcERC4DspQPjRHZ9Q4osksTgVcefbpHBEyOfMWIY
abNLiMdkVxb+qMZ0Jzv+lN8+jJHugNv78ev5IYUhivaRDuJ/4ARhSoD8BwDofvAizsF6IKm6jlNp
K8+W5wBb3C66HU1f7fmucOy3pfT05InSrIffxZ2O/62baxPXBAQ4sW74WtKR3RUsjS6HsCnODUYg
dZeJ3WTcsjMGzAOZj6zTp5xL6lABCR70N9bj0X8dDsrSuSvIRlbqMbL/LnvpwYd3fjtTrwfto/TY
RXQqxml2VA1uAqIvImU+lUqElwqDKKzWDis0XcL1adfOA5Gpfp1hzLmKUpb8BCWPmFG87F+bGzjS
cXOcPWVbFYvMfdeMsJG8oKAyCy7MB4zkMPansRuD1h/UwDTIdPo2FwpiKK9TQc90vpWWh+HNOH19
Rxc/V6dwRyeFfjqtlBRUhcJokem9nMOP6C/sV/2fzLcsjwxJ8Ww9bFZ3X6GhJlJY74gRM6Bx7Yv2
vnbqmK7GqlrwF/kajiciM+2I+R6d2lXS/cgH1xKw1pE4ZLikiNLCFrX6IPiUlPcHP9+wdTdooIck
Zt8smmaW8jggleOjFuz/IinKWQS50qwkndW0uGGymJJ7YQpYYRgSQRTQosUzCm8vCwY8EFwA09zs
63RBnNvx0Byy38q0EyPWCD5/ARYpNmfPHH1lvtNFGJGauUdqxNlJkHx5DFYGpsQpnp6sueOp0fv1
KQGUK/XGdZ+d5BWj0AEyeUKICsCePfn3W6b2ygtTj13KDvjCV1366kR6wOTNeiZ+e1F0XKzOn+oG
W19PIP7AYfKNJeHeUY2a8CpdCgpyh8hbefiuJgr2raCsthJWV5qQlH6YYH2vZglu/a+/ZYP/PYDi
ql+AHapl1YgKI3Be+0fe/61j0qxKZHa8D9dKieBiU6qAnWh0IqwIwu7nfGSufrWwXi6KfuZ4K9M2
0Ine1Y8mDU/HYE+QvXRc3HBeq7uqYWHgiuBOmxVWmQDnD5zV6Po5jehtXlImuuYSgbgKTmzYTme9
HZ16M0rff0KBazEjX78lqNjcb7xMfIRhfqBh7FHDh0RK3y30W5KEPs5HpMEpXS1EdcP8NBRuO6Jh
HnIBX7lN0fq8tqeDFEG6WAEjPOYwo0+39W2OUSxXql1+ZOnxDbcNnagLySMO35vCeDr+ubfTgpHW
GgFfA7fSX6I8Jk64c0ZvhoDK4QQ5zenPS1t1HnRNph/4yywJHIxuzYgFlJ3CGBAj5IMsKgPGA7pu
M5Hvu3kk4rKhwzCz83EsegJgWUPwRbI8JLJeB8AiFekQrpeqXxAodnCOv39u1UelosbmVs5Ky+gB
w8dFGHblz85DMnRWbXzbFkv1Xnw2TXBQhFv3LFUs3mFXqWbtvNXEvKnlr7hSILbADiQ97kgFNnD5
6Cf+0NvaEj7G816B9ID9SN0gsFz3Gsf05y094Nou0fx2dbnoVyvhb2oyYURNEZHHH7VvLzSCQAEH
J5kXUdJ/0n7pUnOcGZlkI78Vqt2i+e2KF1mG5qnxoX1KB8K0FYGSN/nKr3WVW4+LeiZkEfeWGCcR
ftPbtmKV0SqDL6PiZgBTnpbsO93vhOwrm7QVBxhYi3Qg1vEV76FdRXgErKHXDgRuLgsZuRYXLZio
c6gbudMha0QcweXNkTfwknHOy3pDAJ4ItplW3dQ3RJ989MFaohHKjPlq9UcwIgXoysvrRVueXn24
rqyVMJlbxQ5WeedfOSjcbbxVhdD0gu9H9Beg+4ZxLxGVBUUQercKNeBUYshZ1S97C/s7GPG3wpuh
Y6Q21Zu4V8augpRfuXVWadAIZVZ2z9CXYKSj+QflxKNeKPeoOAvqXlR5By7jFPKUksH1qL3jUXai
wZcQY4BR8TliAN9TPBOAvvDtDlqB+cNnsEjH+Pv26WdcxvHLXj5gq60TpGRLCX+nlDQXJweNNGnY
sW5Cmh3sq9jCm6FQi3XEhXwymE5H5xAQj+WMICCiQi8U7AjlcpSp+JOYODqityCKTOr8zK8Z5ULN
ZioduXYnO/RBEWErAD/kN8jUK84pufQJctp1QZg2Ak06EMmh5WEJr+VcsyDANuzvjsiSNYJ7wZTX
OndoR0nsEHdgdPdK4YrVmnVPC2h1vPKg+8gFH5RIVjOaSMfD2Uhgo8qsgy13TAfcRNgl4PhOv/v1
r1IAjc9X4Gi340BUYmueAIZFZuoMIwgnDt0AitXMFbQx6b7HS/iW2ja0ZVAKuFva3dp+3KMPnu4M
dw7EpiG1gES20ZBcJvUPIe3ectMHQPryqXgkcQJ6I+NzrDW9VY4yuT1FvvLs2Ko3O4xp2VLJ9rrJ
UWGKdhAd0fJP/fQaUo+Oo7SN4Vkck+ZfF22SRUySlKaITfhtKqKEboqROdFjvH0iccLK0aBCkBd2
HvT2iEvQwoX/SJ53Xf4Nr5ZEdJhj2wg48r0FA6fTMpw32Fc9wnn6OasF0NIPZ0fSE+N8g6dgwA92
WpSgzTlB6cbaRUNtOW4QWHA8oHJ3tb7B+Rv54+HOpSDnr48Y6/Prbyh0jZCLu+3GjCF7d2Q9AI+K
mV0WDs5o6DImiabqOJygnPdZX3853lUDxI5OrmOKQZoZxgGbL7lPY2NCl8bl/D1zMY+aJ5gL1zhr
yYJRCLXDPVGO+Au70InzLmajKjYc71oGMlid3+Wm/trgTvRIvt/gXzHBxBZDHBrKjujQCRIKp3bz
CyWgVAwW06uaWsGRCZ7pFQcDR0pIoYKNGXrX/royBsMYrfRQz8C3AqqHpV3Zd7BaMYEhADqclYF8
sMfGGrOF93rChDXkCbAaRYlR3kPWC4UvYzyr/wsa0zCDo7D2sgiHw/9YU73X7kazk2B6j9Q61W+p
1grPx2kmNXgLKTkna0MidQ2zxor+EKcNL7TKSHaDDMD0/cZlipQVETscMo66cpEVHroGuaxBHyuE
tp/NCjSz1/gTAm5yqQ9NbhidN9tPzKu3e32Dohv6+RO2r+ff0d7U9/1FASLbaGhVetLxn2DY7WQh
OFJlAskSrFGIZHNLjFw5ZteUhVNQ/rVQg0eN0pwWc8AZ+d5WHN9iUN6GvTV4rVqMBXugf8mbNwX6
qAZyMLbvQXQkBhvPROob56A+F1qna7qqmjW2YaZWFz+nkd8SwktltyESeyKt+0geuKuPMxdlSBk5
WNTYTgkxUtYOYYcqaK0eAADIDsTpHb3TFVTnHuU1ZAmsJbvbjuERONQdEmUH6q3kDXTz6TVdILQy
/nOFMRzM6FZru9n96hZaEHGp6FcAVs167pa2soO9fDRReesRjyjkOk14xdTxyjyyqSykoAZwHN7k
5YsWFlJWfs3gq/BV/h745dYSnLAgg1yPdrkZvdqQzVoL3a0aGpPUd8+UWhgDDE2xqeQnNH7eVeVY
q1NKmexyahVQY0LbSQDDyhHvAj7z0QZc5uf8fE04bcb6TXybWNcGB4OfXRSmreSDc8kyrJ/pdsWT
lYyIRpFemTWPG7Ve4S0XDIDU0DPHrER6MJ9bsivUsjychuP5rs821xXyPfa42QFlbTwM5842heys
aHiPrciHviKoaGiv4sbx416d0vKca5wVZCAU0A7W1BMGMIiCRMdjIgLdDXoULPBq5/imXQQqFj/P
T9VPG+7ksK5U099QFRJHw01gPOXFRHiO5q9uwmtoAqxM/oR8VK5tPbw5aeSTiYQlgX2i7SBlKhLn
NQRsJrKalaMfRIuiMikrNSEqrHCAUGu8HgvnX/4zJOzcnM9LYdyh5vW/C/6jsgNncuJZx6zZwdVN
ie9aqVc32XFdZVBpnWAyQskNdQOtHqj0vDU7joWv9fZz4dQRY1mwHpUpVkhoVtc3fahHAPwzIUwD
PCgMRCzkK7g62QkgwxiGYQRs7VwUxmEelUl948odhCUuvfWUV9wgs/wOhzKguphAND3EyCTvDKTp
0IwEZuKk1BxmoZnvxU0nvMV4JU8mzh817zWtDddjWOvllUvyHuvb/vFbzGZRqdKb3nGfyGqaw2PI
qqCxIUYZLkIbwrk5NI5ucaIMaYyg7zoLE1ZGuqK+7cMawB6cg897wU5FOjTpDtZUUl0VQKqhy8lc
EYk65CqQTcjX+SA63+PUNjqu1XDPN1WbzxS3ixwXDDfL8FqTRbEh/Kb1NRnYgg1eg0VuFNF374er
0gIs2JzMH0+SE7tAwPxuIKOy2PptZ4OS/FJ2RURJQao0o8bQqM4FPUVwszw4Y9dnwPs3z4phN6D4
eAkzW3lQB2G3h0y7hOWvNCXF0zg63rUtCPefHU/HWuMDn0N0cmyttXyRL582+sR0kY0nuoZugi/k
H++Gay8rl8B9ROQHhICsFppINkF9nTE3mogC8FpLZ37Rgat9TSia7d/Xtb+Sq6lFAgBOmLk593l/
xMDIv1o4fsdHZ6Qj38gsB8l4420Gdxh7nUHMa2EczIRf5iG2wxI5oCaCCyiKCt9anat29ztoku0t
pTkto6ByXgsdsCBCPGt17PMS30r7uWEWOdwaATjyb5KAHYKtXsoR+//+gpizIFz8rDCwsDbIFdkX
jJbHYK3r2hXKkxA3B4qxQvR0UXpPV+RVFNN/Nj1D+gsUZLfgixsLS367ibtzh3ZXfkfLzxuloHWR
Yfo5hBo30nnSooIHWy+K2f5EZDCdnLyr6T7C0LCseIZxPuGCXnnGGt9A/eLUwqDEPOb1benEV2+k
qyVn1Li4HD+VikjixlWQOXue/BxZgsqMusY4dYgG1dmYCBU1taiwp+WbpEeN5zVGZG0YgQ/JjTBg
uFanC5J6AERsGqf0LPwV3doJxdnnxy7NEB7Qmw36K1k1xLEWWfF0aVkCXfojkmHPc/kZsKfjT2Qd
ImmpZ3ft132GYWho2WVzyGGtyCKnCCsiFf7vNRPNdheQ880DE41nLA86su7Pm62vOnvHqkXX7taH
2668XQuktxQX4mxBNEOZ5xcJJc9nPLoFw4irb7ERm4wU3oCQZX0aVTkY9oK985u3p1/5plCmCK1b
YbON8ttPbb1pZB/sj11mXULOjRcKNinsQho3ot+TMWAN2GdXeLc3vPf2fSNpq9HmLFS/fV2IxMbq
0B62Eh43r07yhY0ErI4tD2xkeRTet8MezVblUddak1tKH8MiPSE6oc1iQDDobvAZx6xxJkP0AbXk
7jdW4LK61vLMPvBJDxYMuld1w4vBoQq/T86R0ERaL4iSEJRPAB7DY/Nj4mL0J2ujDsfCSAdxr/ia
esAAR4g1mQFKq+knp573FhyxRe4knozXQxD6rsaFcJUiVTJGZqFlAI+Kcta7ggibR9rwwtRhX+Jh
O24YI8qBdlRQETo7D23mGmT5fydmgz+od5lFQXOXqzMkocUW2OGYt+rVSM628Digy6Uv8EVBnj5q
BvBU1NYYlEhPZAHa2DgesXd5jjaITxMKfbp0D8i3nBEhQJIE/xmT9IrkkZS8ffZdyXINuGWfRgbo
Z8TLF3YCiYPDL87P7bjVivLiWgRapI8pYboPzlR8aD1jLjmjdaynDx3qeFqbuqOCOlPCMCbthYnf
rtyIgvS2XY6FG91CWyoisR0vugf4XXf3lq09JejQWfbxEyHyTwscEWfBIOfHbEn4yR3McXf/Jo8H
1KwmtDq7VGCu/G2lwL5jgFqFObdUQT9XKHXiWAgf/72OWq/tEKqIAl0P4U9pDc5P1ZIdmMglHIUl
Uxa11Mvy+WEv5Yi7TkFgyvE8O3bADfqSaDMZVh1EJUxgt2ajupOfV/P5bPWEOE/QS3whZHhUkrL6
D2OYhglSEVaEpxeofNBg7BrqKR/CTwRYCy3WMDebhGwx69lykvfE6VGTRu9kpyOG88vYXziFx8uM
haktGtenYNqknheEGBSGSXBg4XVvhHgGiU4M97zj4kRussvmrHDKJ6GTnXU+tEt95TInBiiSA5jX
Tk3K6j0gr7SzdTG55Ua2H/WvIFAct+aLoBe18rtaYzbOXdI6wSx4diC1ldFenvZM3Xk0fIKUAXyF
jlvy4R4QbRt1pRDj3zPnniq1uXCQVPIgdGQP9ETFBbd2cB95lhxwQNQnza7Zb0/5M4Vle3H/3Nqx
dUM8kMI0JieAZg5vaiHveGkE0MInp1eBX1AEjnJsFEK6OENYusLcYx+6wqdcS/OW8KG60PXxEQvE
VV+c7kTSVOAf919JQqSI5TVO51nDqscfEdrDTIFLPNsTuQ7MXKSTSQDJ5wlO8XdUZv6BaS+sEb+Q
Q4NRNzcU0Ji+VhCXPIUCN/tCSXuQM+SG55wZNPLNFVqhk/zZ5pGC7NGEgZip/Zz5+THUPLRNyVaX
p0AqnfljKKoobrXeNlSGwrLxENWssaJSYeBeC0YBAvoq8Al+Nw9mIRsvAZ1dYhyEsMM8pDCkP6Vd
W931aDID4w5969FHkF54VuSHCzENjLYw36DwPssPTAFClYFb9qXFxg6VXD5lYMjtH6QAzv1fRrIJ
3oUSGEdk0Q94IpxCgcu5l/ptSSggDbDYAuW7yypNgg/w8oWrfJQijRd9ShZjcmZG4rDzAtI6QHp5
pH3Seg5G9c4h3VcF4HAWiiP6AFZBw2xIegcBGo4iFySTEC2ZoUbQU7w0E2uZdSJv29FsrdM5sQez
6o2Fq8p8uCERmktuqnkvkn/puF9/GtyESu0uxDY/KOb5VONgFA2TACD5eiJAslXguYAuRqYTNACk
3DPIqFgGNqFilR932THZcoF4NzSGUAPkemwpuBpYckncR76VV+FPD4LB9UmtMQI/uOAre80evbaU
eK43PP05S6nlD84gNLFPSlPtUM9E/U5ZlPhqWdyX66FcaUYFCyKUXp5kL0u9fFqq1/k0wp2ECRC5
FEFhA+IplNrNa6iTb4gBFyjRZjmR4wVTmNnwTaL+U8mrbXveB1ftdtLQAU71Fx9hjiZv2kDiRekN
VLYr1/olnH35AMs6vhV+4yxP60l4aZMBO0wS0uQrLdcFFJpj2HDFB8dwOBjaUnHvcKBVam27NLWN
tANyOUWAYj29KAUBOFD+NzsPfgPbyF4nKk5+Uq6bN0FfjcGDyrq7sZvhxN9Xyzqr9ofFapRTxTGy
x/mZ8F7K0T+sUioglc2o8EOPHctqbbnMhBrzl2fTHDxgbQ7HNuOUfc3BmDT7yDT/Ni6zXH2wyxeE
zk42v2Mue3tMgc0cannAjZQHxsNHmFzkmUrtxV6BMHjeLj+o0C17v+odb8PL01xB2xGtqMGIAQIH
Gu5vaCWiwNLkonl44/prQ6vPbfvZqDK8Mploubt9/bvHfDoI+Jb8SBWM3/yECVLhr+LlFMoqCMRv
ApBeaXkCvWLqXvUDJ4rGyzI82WzIqcOytRJCbfou+YxOBDz62gPw96rF+TOF5eC9/hpK1btMgTZT
awmbNg8NMjjloDgBuP5lZF0xuo/Htk/hr2kFDROGKWRWnNzumfNCxxVCEuNRicWLCuUABgqT2Z20
LxwDt3s1ED0Y8B1gnpeWJoJW4zHRakNeurYm0x9FTs6y3Zhs6zRc9tudgIqVaeGpuPJ2jhvsNUES
3dI5UD73ob8d48JBntjBk4FdXR/Sn12bkHm4hCF0uVTaJY9lgVfqh/KMLXXoHeyDSZPzBjgyO9fS
NxyHpLDMfwd/p2PrYn2Uh0dCJrnn+fR6QnvsvyldM3HKZRxtWrP10miL8sa31aOsU6ndZiPdxBkw
dX9puU3wIiQyWnI9xc98D2CXckehHDc+WMwiA3bKWT5J0Ue/cpozOP6yzPXe0ZWCVqcTgU/ygbO6
6nYt4s5nRMalYC7AxrMQpzTJXJNTC8o2EG8AzB0R3fLKBZYjENqWC7Ed0EJuGSZeZcpQGD4mzSU1
uZku3F/qI9a3bE/yxitBvkvxZEQ5mWvVfLPKTlaqin0kln/B3f/QyMPAR15WSDvBT5zlDxLYj2lL
X2KEXxrnIpX+cA+PK0kjgh4Mfulf4MhiGHEuIKxxE3rJfEbqF3oRtq/DnR3MRgKvhhKs9RUu9j3z
iPMOlJpVcBQ5xYSevstLbQ4TF3+lV2GMRkepo3oCQUIU60SNYy5BOeTyBPWkdTm/MsNWynUVT0bT
pi8Qi1Dp2jT0JfY+53kPtOIr/qAT+gqdy9Jg6oEzZtRU7zNrfCDcyQpZWmEkqm9rhh1q24fsg/sk
9AmcvYkJoI5xIPQZNLn4D+ZynlmdHyR8mULNrhlnDDiRsR9qFJcH2R/xPLLlgN5Xmi/kcosOChhX
zWPnR3IHJMgEc3NDw1xsqrpRs90XuphylY8TkO/nyn4nojXkTt8bO6mfQ8nCN7/kjGzNazUcRufd
VT9FppKEsxTOXd6enTK32vh6hS7df+ytt4nOto1pQXpfJ/ClsgKogdFSQLp+31KxRODaLXO2hQRt
gXOzQSn0bOKFcp2rswGJBZx1k7RHDkaJ64Xc8FrHU0zCrUB2+vX1NyXZ17mgq4E8X157a0bNkX7w
RhCXbEoq/RWPCI0n5lkcvSPyOc87WGfdDitGT2yxh9ask4ZNi/qA8dFWuZ2M0I5z+PfeZpaldQlz
eOULuaUsig+ZI1Ei5SUAbba8AbXOIUGREEdqoT2zKcIEMNHoXnY0DQGmqt+RVuXVL5gyZVyolgDv
Wrvln3QDH9O8bLWzq6pIAByGo0PB+yty6l+4ra0Hwha7XKYiAB4NKzp2U/ydFrFB17yN1J+kghzn
N5BY3gNjF4xHDcg9ykHP3om8Gc6r9s1u6MfgER2SfSkrAPgxbSAaRNg4IRtzVU1G7H+exAOShZ8y
BUab2cn0Jpb71MQGiOM8hAzuWSdgmGYydgR9Y8SlQUZe2+CK0yxU6F0JbBFU7JLeusc0lrRenwzS
/i4sCCXDWOs56CQaeT4MKprhnozj7ezVEkDE8SCoTGA0gcZXImxiS4oNs/Sn/79pMPvPrZfvTxlJ
sOU7qDwjTosQFMw5BKpPRZPqQRY+854PB9buTrFQabBc0QOxvL+5UxpiKNw44m8rkTHhCeontF6n
KkQHUgqNzzPuiBkG0KurPRQBisDdQrgpr+1+Cx4m/DrvvgDNjF5R3p7BD/l+8x8IGlPt+JIEDZl6
B4ULPaIT2GCM/ewbywn6C8pF+xwKtGAMpL4/a5VapJszdBPBqNIPnRkjTalmSjxkUYm/hDpnVXMc
VZh1sWn7VkpXuL6/t+YmN3WPD6T1DcJ2uAh28CAvhOMwgCdh2eA8IXVdvk/OpXVPkRhREjRSF6Xc
cyoE5nhxI7AOGy6kYbjvXHQJGLbfwV4j7gDKSbTNqU/9o34XzMTGy5BKCVW1HrWXdap2QegGf4px
qFGStrOOERBwKh5XlY7kLBNiDykIra2t6YBSDvO8La7DQm1pJVDEDGNzdFlIRVm/1LJj0jzr778x
LNzZjU06tYinDgmF6VZDMgk0k94c+zwLo+Ol6ocdym5tmjGGuOlDr+9+i70cj3e2NyDsiygxz8Ch
nNKtwF9JIepQ20KlPidmxCyKiIm6n62GYqVytAsMVUvBqUKd9/rWQbpsMBciOKhknIWE9Xf4l9r7
/KzMlWR13RNlmdzMJAC4UJfZrxTUcE4oyLn0PGFr0js0zd0Zii94aD1GGz+o6gG5WlIq4iX9C8vw
Ndm5WYyXwPrasVXhq3a2RKhfKuPrnDmGdLR0VgrQpg+jzh/i+lHTZhO2l3Z2RnTXiKty7433ayhg
53ReU2kFm1LiE5mdXwnh/JrOsljq09J29UHnby8auVt/GITlibNJjPWnLEb5Fbn17PtzKXc6NZde
z51XVq9sEfQzhFVQK3lk6uQsano/b046qunjiCFNJDUGsHp1/kF1mEd8Nn+MB0X/kfuYALTRzKat
pI+cuKtAsRqJ8FE+Sj/tqAicBpF8fjVYMr6wCRasx0apMxpMTp12FeU7JK67VpiVQW8FUPdyEo75
IdD3RyjDNTpi164nlJT4ewXg132/Jzb2MNToEzlsCP2VXvX6YHC8Y0TLKQlBVe9j+3+uWFxNUEej
oDl/MGG/Vn2XBt52mWoJNgWYtKre7SZ8HSl9Aoq5wqCPYT1BDahDiQRxc1tB41PIbvlzK5Uhl9Z2
6WFrva0YpeU1DRrv5hDaZcUZ6lSoSM6EQ/myiTStsQ7J5XnV3gM/6pFKBZjgOFECCesDgD3y3Ulh
YgswHfVeKS9ZZwXzYAlWwroR9Ny4Y6JaDOwJmetHRPNPughDrdnmfMzmDXBlm4F5RknhYrsUR3oi
DGQmQ9p8NCVZknx0IBgb2Occ+oLt/LeJX8Yx5ITHvdZ2/DO2+xSAe4yBM4J17Ey9E0c6NZ8dBEms
r4WNtmNA+dM8SKqbbeJuDHAVwHNbgWmRow9sLvWWQMIkU//DRgtSfVusIQTjKPW3XrffLFSKGmeB
yFUPRdaQO5aWZjtFn9617VFlXN/R8bNC9HkQY03OCNI+ZBEMLRNGkk2kCbG5cJv5Mo698BEcKEDF
1HeTduzY+vWb/Tp1LJvh21gVdYs0fVER3LD1Bg5CJxT6m1x2AIpLTnDohWS0thZPTHsMsyCcLDJ5
a1fW/+O6f+t5+HDRVuuujlwqExnubhhi92jc1+k2k60yBPGkUl+oLQuU3DP/v7bkaUrD/00GG4Tq
I3CZAAyWTxb+WzjJp1OpweqamUkNNOcYk6AW65dWHOzQ7DgFhMX75abNUjun0ngbTxUFsjSVrZHd
j++VKj2PmcF7efMKoUHLDaTFKU42oRuAypFUIJ1kk2bZ/+5OJJ7nmEYq0DFcanOl0Y+junjHF50S
Ijv5B3j+e2CELb74qU4cBfd0TlDMZC4GHNePrA2Fm3ayjUdKtBFHPSiHvZ5nGSpAup4aiykULaoW
mjHpFcSLLfswtiFgkW7dJA9c/pB7TICV6fHc6rbdc+AChwbbyD7PPyWpYitTSWE1EcLJ+xDv1qP6
6oN6AW5JKVCZTrI25Xo7nYgbntps6pUmX+zoOuqQ2IqnoCvZcR/LbI5CDU+3LwWOf7P4i41gTogm
J9pcG4yDr6KCh2kkR7Xl05Gi4KKW8JeoMbmJjgUAlmUSzCBITsLP/CBgfvyuOy9FkoCd2fxB2Aim
lOPKTjfi/gjy0jXajHjQduioC5AdWWwTz7nWt+dtukuI4LG1vMUileRv80oQ2PMLPRlqMyEZBRX6
pGz4a75hdw+dW+yygrwrCvk/T0CDgTOZbZusSZRDxDUc1xT8jEv0JUeZoInXNtxQKHqx8t5FGHsw
P5/rBr2imWA64e5uQmNvSXvKiV767h7B1rQqsehmF5w2nI1xJDXdH3CkDB9+/GBy4RqTl8v+PM+A
x53X+LWWpk9PwYtWtNRqlryxYgK8eGQ0Lo2ZVU4Ag+XeJkY/kObr4YNVcMYgAcJSH2NiZEpB8kkr
srmFvLZgDBm7KE1RsU/A0PiRJKGf5B5YzaSmpEEOcjH1bJ8GE6I8+ZMz8m4uH8JPOEcw0JL5fNcX
yUdSt3ZLDk+k4IuiKdFQ5G1uYntsx+ceHJREYYsF/vkMkVPK5Geex00x3sowJK+A6UdZDBmzzyhT
UqONH7JbHX3HlMQaC+SPciKBgBG81OcyOFV86wj7qAJ7CSVOxxAZ3Z1mwJZAkb06ngfedtyy/P7V
KkWUMplvKZRimI66CA0jvEJtc+yvb8Qjjy1QqtlgeKXXrO2TnbyqPqpqsrjLy2OSCNyuqeInH5Ah
FnOUyTJiD5G9xxq2hoDYz4d459d7urswLDTCulX3ens+YrFLJdE3fAx//cnXQhw/LxilASZkeevD
69DTdV+wP+VDBLJN4GZquqXlMQVUThfzRrWAW3qnQxfqiFpz7oyqfmyeZITSnwZCJeOnMEtsH6K5
fz67xVab1OMJT0XBvN/ySiRk3AwTM1jF6+oTRvsl0Z0iBQ4Hm0Fb2KEyUDnsCCEeUH1HS3owC0Et
ZOqKYUoSc+EaefcY/qMDOGRqdWvsiKthQfmCkvG+vyLQ96NAc3uwX2GjMeoOGAmqEETdBjHYVK3e
Xwv9slTX0psBr8zdhjG2qVOkaPoRG3BQ7oTqVXA25oFG/RlCYyoNxIul7z6VUY5jughM1d3okxX9
sjBe/gc4I/cdDG6dxiVYtHWXlfBn7hwb0GSyT/iAbbuhGjsYmNzMJGtD5Ky2zhf0ta2K8aN+Jlrn
jntjREveeL5FE4YSFjAvASxrzQrft65U59YUsjUT+8ebjXU8dzf+gsTtReT03awk/RrZ8AFhWXfu
epyIBbYRzFwkVmapYVO292buI9o274O2XyDj5YAQJEMB7c6PMqi5r3BtJPj8SlP7kBYIUBP1lfKb
E4FvDt+7DLOdc8acuFofceD5XB2JF+2jyRDPbA1mkEvjkswLH30vSdFtP4qEwT4cPfZJckejrTbL
TvhwpT6FPUYAhgIopaB/F9my6fBeC4alI14+1kgOnfmzQQW1W5uBlC2y43Vq51KX7V837wtf3y7j
PR246vmphnxDxHOFryz3sowSw+ycpSPP3hnzvtEJd+7TDTVyxZNmtZMQylD0QuAMSJkC7q14ppcN
400D0U1NQ1nXgS7JruugGyzIhFv73+kEzouB7UXXv4D0HyWiQYdxt7omJ1TfwCAJutRes8OgyDUY
bMCPV4SHU8Pz6iPgVqnQP58Gq2DCU8hoJfmw/L/bX+SuN2LAFGCRQX4srttQyaqavDJqXMPDsdC9
lsDOBt5oUXpzxy95yNpKsbCz+56JXIArw9f8UyPDRMX3YHK/r/5PZ7wSpU2t5qAA6TVbC507osNH
10EmuYtSVoJ2FMuu6dhhGzoY+OpokLaxRgUtqHAIGY6vf3R5FB/b2A4P8NbFp4FkQthBlvfOuNhq
1/7YjTqxcvTk6746NelcD7ba8sK2T2c3cgLlywfUguedq5LWCrhxs+UomVUk62VdQL2h0SFO41A4
FJ0Fkp0mgLoxTr7gM2JwgqQvqwCRFJXtDPYhBVmzBsd5zXz5TBaGxvp5vw6hFF8XOxDVhs+KKAa3
TWokDG0/CIrHLSkrpZBLfRutLWfG2HjU8EOE65h1qNA26yRQFP2jV95C0icEVTwQfuHUhGN4I2un
IRIQDaTc7XXqMMO5koVpSSSBNxpyDpBgglcJigFx+CVs4A7L1AlWQrrZLNGejr/Od7GKGhZq9Q8a
SmX8r0GQP5+8ncSEmHvbiSLS/G/bxjWYnVmf1vddoehaIIGrTVAoXm3x71hVeM+rBDPGLiypY8Pu
3UHjr5MgsJZv1nzgXhVOL9ga3DeRiWU1G0WODSkGQfFLdERldh0VZJ/FWC/H1LF+Va55IGDOlpoJ
ZiV9PnBgy/ISx0x0YhJdvso6ldOeU/F3hlLpuBBCvQe+cD7k44p1PQ0YYKh9cmccZeZSSyNFTh/s
f2u8wEHybEE4AGjJZvrFW0iHaI/f9YUDycUE5nQTUs5rUdOBAbSFtejsQ2gCDIYZJN2KAJ+7TdSj
N2MkIdbpg2J/4/TMdLu9rnE77h4hYw9er61eUIbVzq9fRn5mR5QpWTwbKQm0qndxVt642ngSZH+a
IynbW+gqiN2hOyVFbENa1LL8BrXyPOVoRkwObc7nTMybErZcMErsfKVI1u4Eu1IY1vyMXuKD+g3R
Rvv2BtYSyYzHVHRvY++zPVT9lcXcxYdEvcpDPTItFbrSPNs9R/QXhzpGyxcfZgADKVJ7+IcJKhsp
ASw9wk636DiA6MRJqJbnhETB2PY1Rz+AiLSJtHzA0IjKQXvLJACktFuZoOJuGL0azNiziwfm3gpr
yDu42/GOUlF88KNtmYsLMIzXeNtv0YyXv+L5oMcBudNJA8PUXm+2dq/CWoYa5LUtUlRC38nh+b24
VDLk2ImTYlmY42SnbXaKIn2EB/9EH3rxqD3A3+h2suQVzmVqi66LjW88qqaYWP8hR3HxWzJyILPi
QGFkoUuDUtpmSns+YjLExdPjoq6olv1zYpHiSgDxRFNsu8StiIhJutCCX/zA9c3QKQR9fyaOYkC8
PLdH5lo7BBKpfo0qL3lBIc8VeQ6vAnBpAeOM6/yDeu39+jWJpA+eks/BPmbXR5ree+gC6y7iiXDe
QaBsaFCQBVyN5eIs8rx0LLlnCSApvQml8P68EgbWrL8uZ2evf+OGpqH0UhuqHvS6H+qEpu1yMjtS
++t15sRHsGzi1mebolPK4NlokXyxUkQvT31jKcNYR8uBWOV7FqP5Yd8W0/Jsgp6FpLCDwV5iyuOt
qYH8lfJdOYmEoN8M4X95c+i6cNE0pql3g9qTfeFI1vJ2NCx46JV+BrJcf6LyDctfx6XEsHp3c027
Gj8jNwqnHsTZC/DPcqyXLr4B55litTHGdyZOlwI67KsLf70wqzMXN3Soh7iToCYGvTogbs8+pJwX
uOMPBojQ0mIaOLC08LnjrBvYLLX9e0c+LXn8A/PU3wniJYMA4MxauewtTCEuDdhI6jJXPuaW1pPE
UwEfjtXtHraCbzZHiC3IP4dOwj/nZ0siQS1zljeEyIirQ+aBh61O6k2VbNGFA1c/oOuND/74Kkdz
ZYndd/N4rB8RPxFqijhOpnaCUphfg4KSVMjj5jbHxqzg8suSsIF6k1gucy16Y82ysEn9lchnpq12
5u7y1P1PZtmFCoVGwrZhN6ARkutmj42vApgBbxaTxU6smgP6/4iuemjxl2js3I7q30xpT5R5d3MD
t3MGoU/lGuPoa7+ryoe+POW/DljqlOqF9l5wBPX5ArlCKo6MYq/xZodF5h9NvYtBGmTSuGs+3NaD
J6S2MNY3tyu7d7o0S3HvbBF2LRKs2hC3xsFVSTU0AREYCFC5LntA0lUgA/nJ9nubHlC6zv+TZ7Em
JlaPzOS2cSC1Pgf4irOAvZC+pGwaQF0QQ6u8iKQUmsHZwJvByGktwHwBIE2jkELtWdBKAfNwcEJo
laH+wTCom659BBXIQxExMr7pYngY6Ii+sLC9/X45kNsOMMLrjcuePverDeu9ucWINyts4Y8M03b7
dvJ00GEcnhl2B39iSkvz0yF6F0q+/sB9zfSB+tL1rTKGKftpaKI+11j6czntLT0aw1fdeDfaM9QU
oQCu8CgIgwdkAVN0tUOetB9e+XTkZrI2fgV7eGjOk+GXHzZH2GptMF1Yu2IxOsu4pPSvz3lIrmAs
ZsG/yJBcRoWW0PsAvvH9iGauPcuIkph4K2fHPNFpoTVzYl7RGGOsZlIze5JsrUDo2Ch+FnJB5ZLb
G56avK9y0DN9wIaI9rvOczppaJ/UV9Hw9rmC2VVLYz1qJMnzCdsZVauK9G8iM01vDGIg9BrR1tKI
kTrDL6WtlhqnSamqUJ/72MUwQKGKXcPwagzvsECAh6bj3Rd14Laqt1zThZUDnu2dNlFwSVD/p5T/
jCu5fi8ojfnPo3/1oLCkZIaXk9Ipf45fVYbyPxNm02Ykx/x7WrZrjYV40iu1aV+kXZXiE1Zd2K5e
GxEA8GD9R1BvA3sD0vLAs5oXbctXYE94s5ziF4QxptE9Tq2NEsVwvPIILYpkdCroeWyIQc5Td8V6
ASxg8DFlvsnLpJAcjAYevQTc6t7r6zfZCP4N4gNPctyc2HyFM6x04W2NCCZJAMP7TYRhkCn54kor
gHCrCiHkAqkhz0nJJlT0qBHYthX2Z00L0YDV9TbrWNixqT4Tta8obW7gH7kLI5Uu0gnzSffPfSHv
B9Av2Ixc+l8gXUMVW6yHCHXL2mT0omi0Ed7OUM2QLlHioMlkaBcSntSGKiDBJSkM1O/oA0Vvloir
AylZupiG6R0kqPMiWlP5P0fylfg0gMluXyb0anAczAbeAE/smrg+EUekAVMABg9ywPdtd6TD13Xk
Q9CFEc6JyNnb9BC5Ur9qFXFGW2FWqGAi/VWY7MUl9A1+M03nYbdYU+O0WWNgnuwTnMMu5JUbYARV
AQZE7yik93vOwEezOxuLCPEa3/J1riftbj9Mcz+Kb5Ays4f5TFs30o6Y9mTNE3PP1ef+6gukhP/8
ABdNq0aOs9rDg/2wPIDL+/pMBTD+EqzL3MKB9LGgOKHt55N/8mBslzR5LXIExVa/OhIndNhiBpsd
/il/SigYd3PCkVkjEtzy+3bmw5GS3eV4np4FYg2mhSvSWDjhic3Z/Wk8wd1y07lagggQ5yHzBN6R
6LIHRJlqdpn/uohlfeUGgs6JeCqiPv+zG5joGsc2gUBPTlt0koJAByII1/0L40HY6gfH3BZMPatA
DEjZEp+M/Nom2JupoeJVxu+yWMckvD4QFmGSfYDMPZGxTQsD63A35yBPGGpJCvXoc9dyFqkPAKsz
1Aov/Xa180XDrBheQifyIHxsytzjcYCy4QmZf0dMpGCyZRKtRbsaDuC0glvdCmeS0vGHSu5xkuby
Bl46cylQGx2sQipGrVVndF56fWQ6H2I76sxyG3MdYEMa99GABd+qRQurg9P/ch5FbW+SIKrR1kzW
w9EA5LJS+G6JdFm9WPa2Mh1hd3EhzTC7C2qLwt1zUTevdkSctpZbeqCe//Gup7WmL7BBhUq8ioPp
aNBFXp7wBSuPE+yOeLSrXm5+Zyuc14vVZXfj7C15J0stx5XH6n1IznEWQPDHZKyBphOy9AMERNle
T5N2rTm1n2HQj/yTZoRmpTS361GdC8QWgNA5Ob/iMoqEqcCh7e0VGvwvQaIi443XVH4hmQGgOMuU
vDifD5aFxa3o+aF1ixZNGkdq+0geZPWsBTOaqfRJMquG2mrojK+mPoBRBFPLSJv8vvfqxKrSkWUK
9CT0ynxy+Ehh8zcTFhgy8Jj5rZ2FCxRDFi9TIjwO2zzWkwuokeLn6Fs8FDQaVcOXEPVLSNYw8oWh
S4P3/V9ayq8WuvbotfNtQVuiwJqsqf3w5NbbCZUa6exgyEwlLBK6ov1ArpVW99y1J8tC7fhH/JJx
E9TsniOmNbSbudYR5D2XHF5qOyb4akhpNKtcKRQ50TXXQRm7gNVdeSrvCcokbNUSiZK739y+1Xmf
73A+voz1WGX7dNss/ntGQWmMo94nwozhQt7oTgmwU97EzFHX6UicAUgF1HEcchMZcOMkFd1E+K9F
9WLnZFzVlkDTR1b40POdNysLymEU0zfNnAvTqHAtSqRRJhboZOnzxsz42Oy3fvJqErdtuQpq3TJ0
87dPpjhPAMRFjCZ+NDh33tnhwWXahvW3Ilre5+r1VBb7wsnLqF8kX7RSGwaRgzQkpieEXcL9XghZ
YntSU7DUDci66eg/Eb/KbkNZ/9LIkw/j5k9l9vZtenCRdElYDYpzszor4F6w978po8p8sYNNSc+3
XIH758R0JNWM9VWFZS/JP89GwuR+Jcq2n+HKP3YKukGUC/p4QD7VYLlzpX15mZ1yMFWvN6EeMQ+9
U0tjoxE365+pn9yIa89ZmjClqS2xysaQi+Fwraufm5ZPKCoW3sMMQU1xcVtOIFqrwQJEUCm3mbD8
R+aE7kbAy/unbkE6YgT0HJWeVuJuFhe1O1XUHiLlUAEgLDsyUrhAhqjBsQzVBcXorODoZDr6UWbb
yD1+o/60onlxCBwUtkTw++tb0aHgYHULzXSx/CfRGTqXBZne7Ir/XuElPkx+sobASisKw+hoJ5HT
f9eLrxCtJYGLsb2fxRZiREhf9WaD2+AmsJIMtEYYby+Rx3n2GAwpw3XkJTCpBGRX5j3yUWQ4sLq3
ZUQkRg5zRwthKb8BkHf3AcM9QFQY6nn9QWCiqKV3RKk+koafN1RRriHDO3ZzGT93qEe4676/b0CM
alq3oLzoXhuAW4M8q3E4+oqnB3Zp3ka/wp3Z5rarYFapV547Kn8L1keCzt6Jn8h1r9jdMH/hfFLh
zpuwns5zK8PjtxUaijvgLYszeeCtqusKTreiHEj/H1kikx6XEhrKV7xg915gZ0/rBILzGaIFiDYw
Bt68ERYLaPtQ7X+KUKPHW1w1L9LJynKekZD/KHs8mHT/bwyGhI0q7QX2rDCn8VJ86OQyO38cR7lh
g9A5COWniXW75bJbeVf4DXxh/hODKWaUJoz09gB8hBxmeq9iorh6UEYMjd/ACGPQTUGDweOC4d7s
t0jf9+PFUdC4aC+i4UUVteVcxZGOgKmdaNVFoKR62DzqdXP6bOamkDRPAwghcZNca2U605ay/lFd
u4d3Vpm3iWx7STcnVzEGtrap/2BR3hbQZVsmzP1VA6g2oXAnKW3OsMbfWhKGE2MTWguiuI2EZRs6
b4cbqjaLwnA21uEummVHLk0tHup1gFSDZqGI9EMNWbGG8L4y4yTYAcncwKzli1AtmsaAJZIB3bAQ
ggCn8PJx1DaHDw9g8zPs7gmJw2gWftIUvWr1gh3Xr7MIYOrr05OqEBf7ymSMTXhLiw9ewDXYosFh
rHxopIjHKBDgwwYuUP5pOZ8wgQFfemHI1gWk7WIJ4d3RAa8H6l4U9/IzjTx68O6HKGdlnmPc+a3/
elvZyLbmWCUR4qBMUY5jH+ntaJl9/9WWk53EN3OlnBfNj9kfDa6zUTRDd7B4RniI3dUhrSOSAhEE
DwagOpLmhZGSiTodhQiQ0mBWMs8LaThFLrh75ZbP1GL0iWU/l4NROqQFr0axMIdGDMw+qTYb/iIP
EzLUB2YJQwvhyVDViH84Vs0bAzPWP2Lq28/xQp/4u89UQ1K8QY7wRxeivlkfjnHS4KegNOZuUWFb
umeV+QPcOgO0UWgnjgdht9MhFcLESFRRqSWK0HWtDxqcQjfCTQaw/9wbdK7z/YrbobNyLl44vzI7
3HsAgsA08TFMvg3iZIplYDhbpYW0offC083Llgmpd9pQaq+SKDtmL/19BUdDgyiRYmdc9sl/qRaR
/qlC+BbYl9fcYY3VfPQrvv8lVGBY0KKqhl5D99xWLy/vZjlZ8qE/DJ3/q+ixroQEgOAoyc44A/OA
ZDS96XHk5dSIUUOjUL/asQiTmY3pxn71dtdOp+aHD9B/UGgqRxvGwypFYokhVMeVL2CgvvRie3tS
FyTQAMsEEL7PbuwLh+gEfNHaEsAUb173SsdWAG+15pnXzPe0CQ5bJv9nL5LeuA5U3mzaOFDxeO0w
ZrKLjogmbvQqgr/83ocPw8RSDxui7IfY5HKpGQiamwMrW16WwqHGxLT92N2/seIVhaqcOhiwCcoD
HxlAP3RMjuMbaJZeWcaxdiy0USxFGCSLuwXMXgRyxeHWu1FciJr0aFWgcrkWQV6EEBIRq05uNVX7
odmN2OMgSxZ0zJErHszRnxrrEuQwvLGfJaRDuFy9cHQy5ZM46/4jqJ9So53GYrdJyIq23O2CrtMw
IizGCBqF5oEa5fZu67jxDcbAdpov0NbN+d1vFUJgLs19Mf0mdJKN5jvpzmwFJ1ofepHdB3YPc/at
V2LgBDAp/ZowxlDxnul+TbUxUzUBeUlrZnRvotwvarz/5nlvaM3AUuizb4xCe0kLJjxEEMCMpJ4l
C9LPaLIrinmEEpRcyTz87utDOOXDCSrBFfh6FJLVQ+khft8bjs6UyFUK3RjBuzDMV8JQRUOGdFSR
pJmDRT8Y1BVuqQ1pxwCAWoW0KF9YlzexHL7BpyW1dqfxkaDOU9kb8sufhDe/tbg9lHw7v6zM5Puj
t+1irsiOhf4sOSeUWjmdjsJ3NGELUaUFIvdSVRmdOP7apAfwqWnHeYLWWLJXzrGkTmT5d5svA14n
Qb8BgqsvfPwOmVPEO8obRTbAIUkjSnrcG0kVXG8LmbzYNa4zWeg8j4L1K33peNiJyOKHLdVDdu3O
vuJlth2s193qVNEbnGn5jEFTKtSCByFIOS3eGZDF1vT1tn15FK+RQtnS3IKgQgwfO7eq65k3GqxQ
5c/gC8pyYtn6RpEKT5mCCqijKtV5b+QnpS76rw4wobBVhTx/yWZtWudWsAS6alxHgbjpJhVe0ZQS
8Tm/Zv5dJNCifmq75uR/sHoGWDSbxYrrT/GQwSC71UTLjVpjNaJK9W33BAWil0IuPoo1/QH2YrtK
WnrRaHVWLkvKe/87xEKhENvEv8d1CW3lp8qZ2btdlnVaWFXRk/puTy6YN2siOBCltWQVU0mVxtKh
m6Mp8rEiflP+q4Vm550aH/HN4XcBFAVMvFWkrk8CHvnidxRjNFkXK1n1Rfi/CeipCBIklA14SfaZ
0R37JBldxVbbsOt/RBjeWKvcoSDMrqIlK/8PApaLjHcKg992jv5YJFg6guK7JAnzF61W6ohmv4eb
SHze7qSvFqGOBiMUai0QtL3bzscZCUcd8fc4emdk2g7/gj/vftda+r1kScDea0tKG8RuCoAVyoxj
JdlRprngAIHkKZq0xdK7zbtRROZ3KmwxqeSb6lQtSb3vcWBZnNsHFCi8ENh/7D4r56gStGff3aaJ
gdxLqvYD9a/QjSe/qz4IFJxhVV832y5ef4ioswLQeDE+TxiGGdIuD8cjKukp10tAax1P5FfUH/6p
Q7vAI3fWy2eBlxZobLuyOP1JeF0mjHy1KJRn2amTXLmGlKtCypHBtYdb2p1is1X7riU16DDRxnAm
az6FD5PoQhDMIh0XlLOrjOBfU/sDJAukB/apD0kM4StDrpv2cYpuwT8aagnoEjO1jitTU/jMUKJ+
azErY/mld01Uyvh1eTtdlcZnpq2Y3MGswJfYWVAxQtyFa50R4su0oz+AkGy/mg6aDy3jwqjPno61
e4tWUGAkvOOlv1/jupM6UbQ6USCLpOhy7OY/vkTmH88BmljUYgXjwUvvoYRjxfrS/+IvwLMGI6F4
LsF+30PCnDryytTYENxnGo+7nRnhJZhuoCz9GAKOcjz5AtRnfIS1iU2r9+1JDdH2lXR6WMqgV73k
KwNBaAfvpJ7QnuLyDICBVwMO2+mfQn0/a8m7+YRSq5vz8KWYUQPHv7S3CDUxIe4DH862T/taUJOe
Tp3E5G/OBpHhQn//tfMkymsn8pDMdKFKtqO2ceHmG71le3DgVSWMu16ry7D3KsS23RRZ9YsQkl4s
YhX7d7I20lkAQa3nWxGNHwMtZJRJhM6kwTgPfa6Kn55tO3Qg6sj4O52Me77zvKY3NzRw6igDg+BU
9cd8pHz/MAHPqjS/hK0m6NzSDtKjc3JRZlgGutD2ysZtTp+ynf5LG70S2+4Er9RSYuAFRqJXOp9T
CR68ZhfS4ksluFESvKtdyxpEbW/DkJeGuy7TTtGl4mH+pNi0Xa2kXg+280DoKFedBRkTFr3Cxs5l
Tn6dg0jdkL2kySvwu1ELJOMn8qjxiQs8ouYEt9Mxu1qHrMsLiKUHpVHWV+GB9SVxKalkQWfLbjqq
385+vCuSoXizmNqoUhCPILNeP1K42OzIB8YXrB5Wg3MJOE+PLJ3sWO92J8WfExVzEI+I5jM6z4LK
4w/uC/huc4v1wwL1jUyiLDiuKu61GOS5EHeAHQB5ux7LpIRfaCtY2MwiP9zHX/BNSwVyO2FbxLsK
gilvheSiEE3NYNl5qDDkhW4A05acr6oJVrohtob14CtKyjJPfdMINZoYj9i9G4EG1kU0DPhKq3ta
8XH05bRDOQUl57ARsQfALrEFAFYL1dbRJnYirGjwHVoOxGFTHXIC3eLHzWx+1uroYwY3IdyJXWnT
3xdXsd9GfBGqjR69m+IWQAcksl6jr7FowzU2acRviam19MDy2gllgROCXUHygIhoM9FwNrHkTjTH
FvZGp9hQWXceFp0yZV81AsMvGQye7PMjRs226UL7N3A2/YlikVVLKUkKzPgAGt0L2ArW/Q5tHo/2
m4+y1zWghbZTIvXN1qw+L0N9CJ0H8l9Csa6wa5CJpXbJstFR+ogvkXdI6lANHkAnoHxlM0rELhiP
AdcAogCvJxE8EVUpivCSCQDrZqMLTpCI12asS+u3p2X6hfWq8NfJj1nbvqbXRabI0bMoZmr+YZ04
eDi1Mt4lDevHgSYst80XWoHCW3k2BwuWa8FPL7fkiz+bbfrF7IElTpWMH4AFCibg7q3W5rnOUl8H
x/Xa2E3L/WXrumZVQl+jsnLxDoVqOnE4lPQPxyhNW6tAMk5QZl+I93AgYSL9kG5bpE6dQScH4eJU
B9NPpwe8u2s9CW/YuhnPHdHncgHUiYt6V6MfkStUN607vJMw1oukMbWc8Sb0CPveYhy14SXD47Ct
BaVHahJFNDPmzJrHH8tRz7Ph3CRUwQ4biy6WfokpCqBfgkRURnF1ALto/mrv9VU60bn/NIzRqdts
f2abPUqCaUAsyWflw5QotKCYYO0Hlbw0hEhRTfF87gsm39fCf9XJiSXiaa7qzR17ravMnb3UE4Da
7VytkGdlXdqq+IcJRriwZaxgm/ry/vt2Ez9Yb6CBPY9/xNYRAm9pj8TooVvRXRCDcgqaZ9vEIazn
mS6ceRUU2RqJhYHLu/mwjMpNBfNi/LuZlR/L85AWzeFBjyBzzIddy2qiITObZnhcTWU6/5Z/DSY+
uFd4O0yEkyEpCzjwk0Ybb+z94Ow+pcNuPSdJzopUB1uHBtSTj7lvNP/AwAx/SNfX6gyWvSXxcyfO
2RResTlwsA3HfN8B28bmeWdOqXWiyTdgkIS+xce+FW98+EV4hKpkNOhXjcvKBv8FdFjIZNgfd7xb
cEM4GTXS2+Mk89koMiNx9ytYKftes76MQMz+bmWUhZQeoaa5iSH2FMQ7QibVHG2Em6WeWy9iDu1u
fszZjKqzMIdBqveonvF2SUlczTGHeAFY9B9djTKMLkPiRy8Pfm0cUIMdA8fdX5ZIkHyv8ACXU8ip
sIYbZj2eQmxvdksIfPSInbX5tIhJDRFXF/HS93Ni3WzyOQFWGytx1TNsYkJMQwlxM8aho08leeTK
lX8zszT6ENu0Ke622UJ8mQR7BWhCIKK0j+Xl+OLSrtU9gC0WuEJ1pJrye+1ArzbIub3Bv5qMTnzi
wgRH97JtN8nTDy5rdcnYtr2aKhdSQq20gXVVqb26pdK+Nj21eE8Lw0/wXr0dKPDo6QDoUvjnvPR3
eNAbvf+L39pjTViC49gT4X4Ky9CmS8h1uR/UBTOg9G0RFL/ELyW6Ht/MWb9vXgrAu4EgVwKgO605
GnuuBof4lJAeMHtikoowows/BHGZ/l+GSri8FndGPza3c25rJg5MBSXWSw4QRw4ms3/Tl8oyZH2o
SD4Ob3o5fYEiyl8njr8z21jnXUrALB6La5eEbU5l5ImRn4Eiu13BtCR8TzIOcMSKsbejKwtlqs/l
Hm3j4d+tyFAgyWTCqOh5p5ojW7KySOKfsl9fJ3MlsmVgM2WxwQufF7IDEdpzdxdhtP6qhUkHsNFS
MITuQO3DMh0G7Q51HNa6LHJXCfJDVAn1cut4eicgTVCwq77TROVSWFoCbQWwC47M/q6ZykbtT3WZ
bQsSlrUjiWEAX7ZM5VV/XO7rB0tZaOLwer6JPVtheQ+Bp2Sq+KmnFRjZAheAzHpajSTqlW2s+nzE
cyPzlWf6565sPXrjjRwk3iJSdBbiz40NABZCXFV0IXaCzGfANz0nlVBnpMu9fpdSGTkzFbqOnYXm
FK09P5OB5/yxAeWOSID4o4QGfWriaa5RIYDfsPxbrKGkaRudli6/E04/haT6WcQO1A9ziU4GdvAs
xjMy4px5ETCWxiyxRKt/VM8NzPcsisdi8a0BPq8JdUWy6yxVlVliti959NumW/vmu8qP7R45VV1V
jpaEW6Xww8wUllgLjA81RQEVX1Z0u2MF2gj/GNytsADGJ+y1IBmdv9qfe9/eKTdNxTEpAG9+1FuQ
se7oi50PkUYwHSEmAWJKs2MFDKev9/Dhi4gSUEvRKThCH8nIKELAnjONahJ748AFGtu48YBe6ote
FEIDEURmET74rSCLj2MFdg8fT31FP6m6DImkyDXKRiXegxbxK2p17Qg63AyJ6D15CHBpxEzxm90a
c7gnQvZrGUls+Re3W6oDE4O1pql0/xMBvcsetlepE5tevJRdt+4PFdJm5uCBS/qF/+ByH8Y3UBNs
XEN5ROmhbuH0eCeAtB3eijiAJ/KgKsBCLLa4Sl+79fyfmyNVPNuDEDP54NG+bKBl77CrAxoOXw9m
ZBm78nNtYdlHA5EScPcdS2UK6wk/jKf2sCRmyFqM7+Ttvov5zlb/Gun4bUcIQ+HfBPjJXGdML+AM
+tULbwNc4rxqXXoseTD6ecmImcbtLgmfsrT6GHuFZS2PWf4rwrW1hmAnSKOtcoYTfDbOiTpRfihy
ckKNDvWjSL5KHuEtWUx48sso7YKjrsJhWlr6Fnir8qs5i2cD5QQ/0GbUPggj4UEFp9PpuiXHid7W
+xaCuRaajuinIknABCq0Yu5mLHiW0eyemVxfiPdcv7rx9Or73mz4J2cWY/6QWEnhcS4ZJzPPWJUB
+dB+lEipu4UXM1shRZoLXj7vsKFff3MTcvPQHwPblEzpMEkt4lEbL604f5xVhx3j+TunOvwS7pGP
RRwXLrs7qhjNWsMdh/CQ7I2/76k3DSS6k4zFwCVvajH92DdAW4O09ccupdWT6fx4nGf+DLhN5cXA
YWNJpK/hIMoAyDrI1LHCFUPxZVH/wEusJymY1lIp57b+SEg65/mlfxLOf0Yzv6O2vmO1aDhMFCug
vecwaoh1mFvSPbFb8IiUwI2hGdelGxkDXOBkN/IZGrdARV5v7XDmbxf5wFiDtx5Vj6hWrlPF7aoF
9GohLzUNkVvNOCBuj8DH+c21R8mUS9eWLFfRQekCvorFAlWdGlrkxM6zI6vDxE2lvo65qHIlBSUr
Ahy/3VJPkgfuHlT2NG7qwghYyP6KFL5UhufFUSrT91DsXjtfw4rERMDF4t57OsYXHDo59/fX77Ie
0JiuOQ/mHdq46/Hjla8DTI9KHfB03b5bAYir3VMhEl9GaNKliXC2hiUXCrrh9Lnitj8HCxJTvXvG
pUdTaHUHxLfxG2hmRXQBWd6LzbZOzAdMJKPuYWK5ODWO7FhreyRGiTEg187CMW0XchUxRaM1A6Km
5qJBqeSFGKmuXOjBwDr1xOY/4wDOAXbYTdWdO/Gn0Z+8bfOSmxQDR6Xrbrll6/efNhNPwvjDKTI/
pL0XSK0waiymvoNLhPad5aCAo1+gA7f0JQ4WEcMKD88iDQR3x/Dx3ufc6kwGA7J9F3f/ewVGbYKe
fL9d6/bL6gCKcqiwt5T67dIb4WcCWe70gNQvN3xYZhXwkeNhS1x6uVPkg4EX1VR6XLcFpNyUpj2o
3OaM0aq3gt2IuuE/kfIenRIQaIhFyJTNU5y+j+D6anRblVIqLnfxjxWb6POGVzrqRTIr6K26oE/Q
v6jF4n/htZi2BcRjnNbb5U8OqhfvEOA+3yDJk+dM+PAfBbbgne0vDxhjHZm2Mk3MtFeo1zIpHs/K
s0cVk6Ov2/fCICXWZrv7OJTH2BBD/9H1nrRXT114k463dzlD+kBXHqycjtz0XLSmHcpDY4MVm2aX
X8Bt+SZ+qLA165Cs3caTQJk5XHYsrOQ0yevChvfl6aMQsuQR/sAK7zMst3zz5VhWpiC9FxCtidMC
KpEpXON1GE4+9+qjTRc5jF8VRowj3bjrEkC/MT+jH0PwRJfZxiiFxfO2A0OirbAkwA738Haw4fOW
kRBZCyzGJ2YM8gVRIVvJCxs8YqmJHI2Aj9Xf//95y6CKWWPGt1H6/8y4lBfocf83M4r50nN317mq
AIlrtkH5fzQt+TemymvuekFIap3HKUTxgvllIN89NbP7xmiufADomfRFhuc0lqSwjMGTpWW7i7mM
2F2Fm14AtOip4UIPuZQylXAIrcL22KtpvA3it35nFEKAAwjI0mejgtN1FcyRWhk91CD8yEvWf+v8
GfDuOKYploN+SAq+lVWkSzAVBEr6VojF7J7SY+T8pIMDrNOXNg5mxm9TYm0/g6566IbRjY+2mtm4
uAl+yURO6AOn1yLqtnotTAntDIHn0t8tHzVS+txRxd9oLWVFuMlDSWRC/e5EzkkJl/KVR3enBGyN
/3Nl5eX6muVXZcCaZeqS+EuZEz8dWQ2RQII/UNahRiMTEvP0TJcLnCuuUXes4GyS0rNOr2skj+TD
9/0SwFJGwg6aEt/BGwW9LR95d1Ta/+dQmlo3wAXz0cWN8kbjBsgnUgPYLZxQWWKlXv6iqD2z/5x6
0t9XHGpmrlarLdJuUSyxNnBDx5VFZ2LWDVaoe6r9k6odnE6Gg11oeDwyfkPHuCXXJoI9oKwzw0By
MP290IUCdvxCSJtH/EQrXfhl88D0R2JDQTP6fX2cS0QnLYrPTCmrRDYEb/E4A3GHroVOXrfu1FJq
bmI+73bH491Nnil5GyJOBbFNeE4RwIkuJ/me+i/x1nB8qXETSRctoGKyPS6Tngln4qr/k9Lf1Gk6
UFTkeqec+sIdl8UosIADiGDt8w1mTuwyK+iiFznl9D4v+rsoAf0BQtl0GCrS6JKH30WuWpVsmXsx
EgYaTNtnOdsNMMUlyhhSoc77+PtEiAxK3L34c7sgNmCVprTaRS6Wul0iJBhSGi5t3CBOz/1rnYvL
oqgy1kA06laqIcgaUM5+R6Lx3H+W0gF8LZIl8SbiH8zbMoP2BTx7WNZshuABx9u7geZj9j+WQJ/O
mdPjDMp1HM+L0/QW081ycXw2LG1f3T7/wQp+F/ng3l20+Eg+Yp5EtAYQEEJgfGFhOdSDiqnhabfE
R7jNekbeNne/tT3SCoxkbMIX0fhAAxVO6Py7CAfCUHHtODRVCjS2b52J8vsMP1xiuhEokyBt0FHk
NpVHD4bS6zP0UvIJsbhRFzv6/+sN+3i3RxrQWMW+YxnBJqGs5y2UjQKYSw6Y9LEvKYJKrABSiZkL
mqCoVvbqLBTnXa/ZlqkVj9O/1DX3OlQcKzVg7ZB01PWpEjeMd1kU9gbPAC6norpAdoGyeK4aa4G7
Vb+5a0ruavpNGIioGcu8p3z9RUGIdMd76HyTHHLZh4NaQajBLyh3Qe4z/xrGIjFKaOYVs9fl0WvR
s5V9UtUsBaZbnNG/QI84BYNBN6jzH+dWhXGwPO34g/CKTwV8840revsRH0peCJdrfNKRQK2o9iXl
aFnkx9HTYhfAN5LIpLLkuQUZn2r/+mSC3+smwHsmlAJP20E/bjqyou0izLHykcehUYFd0aSHqldr
RnDQrD3I5p/iA2qZqUHndaz8X31N+yO4GrI2N+z71OtICJg7ard6WtnT8vr9wDBet0AlNUVY3cKX
Uv5vE7jK1FYVQh1wXkbstQdQ8NJTayT/iYFz4sQ3jR4iHpy4x+whkVKhA8dhZoZljrpXiSpgrI+p
OUI4ALO2gtUi97NobZFaPBohUDWBUBKE+92ueHSxLxHkKSuk13rM2VbclvXBu3151vG5wOq+oBFK
TXkdjtjga0+zKIOnB3KFEg1YJN/f1TKBgnaS3+Y9oJNQ8ZzOxF340/Gdk7QPIyBDnE6gm2gOEqZa
VdSq/FcmbR50bm6ze8YKb3blBKbjvhhwsgDn4UCCHKMH3P0CncMMSmYIYmB19+vnYSyI4vu9z82Q
q3ZLS2uXb89hyIuiIFVHHfRVVfzn2JSqdTJx9AjAx8iixoxVcL++DgT2kvr0Dh6jjANStHPYmZWy
C1Zr8hcXkezgwGcRhVvLdiUbEuzLryQGsISYQffYTjalAaCl0pGzizMhR01x/uKe9QSS8K0NuwTq
wAVnZRKhuuHQ8hUYnVLOsfYvglp8SYsnZ1tjVRH0eN6NUtzu+IjvTEOC8krl+A6QIcv0PP7xJ5tc
WMIrzqTkOmp4ly85t/gUnSw+MNSrP568QCVRt5ytA69j6bHMPc3FyHTg4sRbrS9zFDX00hbzau6P
XjrtvtXru0r9w1rRBPo/DFqs3NuswJXWgZ5DRjDxR/T50FVEUwxME1KGNV9MHb+FeG6zyvvgQECO
6sQObkGnYLNnwMtedZgJWapWxbiUVQvhDNns57tPvhY3OS43nyKIYLj9XfHn7pAN2XAjl2cHKwCk
69R7fUcoMxMahMjDDeYJjdod2eq6WxPGoLTLGYjP+bsWJlwYIcEZAcLmmpsXibt99DJ6A82vKEyd
vpY4QXMu8fsb3wzIDs7RoRFcy8Bpf/y+p4x9I3dwWsqUf5YoZ9aK/DkBbFSY1neei6vGKnkfowVI
mKziKklISoajfo1Kc+qzl8P5hM+afdYKRS8DAi988oPNoNy7t9c1UI3dMPSaYqK3JgYWo1B9hMi+
UuUbuTa0M2JvwjzPu48oT8RAjStM9OyWexZPR8TIDu3GI4Goh4Dj0buvj1LSxGqE24EFpGI45bmA
nZjdpa0s2oU6GzkyTSiDKcLE9c+tYGpkuMy9O9A4/BpM92hjo/rxrPJiZFFNFtAWcsTRhqKirFee
fZtaj9XcMEaUSf3f6zQK2Vj6kOcI3RjAiJsuYeORQDa3vuhFfOzzJN7goJr1RmAZUPHBvXGz3jrR
Wwdq6jWDnISZTWmXB3GdsCOXDlH1ixYP8aVaqPgI+Ky+eVsOsZQK1LyK6Y1CHWhUn+6cl8KdxKzI
dlrtRUztCXgnzPlbjYuGnnguMYu32k2lN8pwbXQRaLOHO64tEb+ejV9lj5tQZkSP+/x+swwGbO2j
FY7qONkxFxTYliWBuWCnNJwdPp01xlTWaiYdEy4J3N1ZE1khjxVmMGJ0NJL34bZAjlBFYxzB+Jls
c1mu1FYGxaaa+f26nQwlbwY+OcfGfDk25RJPVoKZ/VUq9Vb1WXWln7qujqHY0S7QHTypHMowsA7d
nl8FT4nuSj5IX/aClGMPTpbS+z7K3LSDyKgkAM+ooNAmZyWQij0QJJQwqHSXHXIrg/2DfwXgTvOq
EA+fdHdTh+zg0LggCa/LYnBUO5H/oAiC7scWdmx3oNX3hetVDafyzK3bVJCYH0lcxkRNHzrs8VyL
kxeoCCLuw6O16q/Fo9pSBSgY3k641NJv759rb2y/OHASluEcyMvID/lO7OergcVfOseYdG2rviyB
I/1RjsNWzQ2HY3pAtOvWB4t1ZlArE6n/zDctAl5sAjfcAufwgmmbcwvRpqhDZuY3tgcT25mVNSet
kf+fOBS0gpRhpzhdzF95351O9szc3Sqaj5bbbcArKRWNl1cSk11LywoRd3RMGlNNny4Ew3jnRLJf
6XcKFfJKARgcV1yaAB37b48rdAfcuJDyGoHmpZLT1ApXPi6Cc845Dh5I3/G0njf17/VYydtxzagT
SrVK8hlAS1r8auvMdkQ66Nj8xbrDgzzA4NbsSsy+4RMWYg8R7z0CHbbXRqRhiyAR2Z8i1kNbWgff
bM7pUwmxvxp2Q2gGDRi+z79M+TMLlTl+s/CNHkju7tleBJgyIAl09rSue2T6qFkrQdYwFj8IUa3y
ko3A7YeSVqYuYySop2LbFOb0lAr8RnQ6EhEgCWqADanyv9XxnGp+gIDY+LZ3mCx9cfFaQWLRyGkb
Qxc4PLZMbv9SRPcMhDVxVAFtAt6wH6EpogPTEhmdf+PIZ0h++PJNNp0OQLKkxQ5SxVILqrvScWk4
u/uCUGLZ8zeYhfXmeqegnsONmp1RLoEV/j/BKARaTsZkHt3K69CceVPTSsLmDn7AtshxAs0yb5FX
zuESFRHtqH5bpXX42WxR8a2iEyFArdlInVuvzVH+rqiMx6LSkqVspU2eadl8uH2tn/Uy79ahtfPq
bOpXbMsAcXiHbcQB8M/F2Uxkd0sD2fUmq4vCn4ml1ZevLnknblVfRxyfEG5s1cPhmrl7CuF19EwI
UH3CAG8tuoBec+NX1Mh+LTAaUPS7oJJAOVOVL942zhPf5ms4f/MiB3q6CyoEjvUSfovAsgWZQTnU
VHGZnwD4n7GdJg35UU3akIZ0kVFmcSEk70lEEEQ4sfYwMte07SS1I9vwZ+LSQzMK+V0ztTdZ/Yf3
qNc1BkHrTXND3cEMBkBfPJ9AEt941RtRbBQvNAHk5am+dCecbDWbByPl15OpqoTkDjmbcL/AFZFQ
WhTjK4xkf0rPVZSC0b87a336fIvHnIaz5bV36zxonRI1jQbmlI4fEwouMIbK5DcOD1sElTzD65KJ
EYmuCOgwrdnnH4Tc+j4yh7kgTacmRw7n128V05I7aF4Sl5Kw6aTKYVH2gc0V0WBHFX8ldsUxZWAq
vJhLx1Gexnu2jJO9CeL1HcgYZbGthZbCw64KKZo///utiaoEzztlkTbVb45n9ujnFhQ0Lh4Jx/zp
T7U/JvR7ilfU7oQZk2ubxHDp4E6r80DsAbC/VPiSMSL2KVSRA4fXJQcIkxxRf0xzzKTMwrHd00WY
Oew/3xdBGubHz5XmZ5zoLv+wuBb/GvaYvVi5oS+EO5Yn75VQRSnw1GMBBLFtmErrvvGJ0DiQ5iCL
Xit0S3GaussYshqlbRSmZzg3/ZbsW99q8dtyuALh9dCDLHCREqki/ZdUEn9zlRy4obBlvpP1/4JA
3fGj71ZoS1Ae/TxyXiLmhl7sCmt6jKBbMPSp1qk3gLLCw2u1xbLuVMlGHXayuAI13mg0VG/d4HTz
WASlmPXxGzeWm3oauodykg4uOQbxGVGNJbrm/rRv0liPQe+39zzrd8vCUoqtCnVywaSvUZYeUWd+
IMM8H10IrtKnz8zubG4Gu8MVO2ygYvaKaSTN+RXZyQqKyYrABxjWFwjUrn13spyLCkucuQCEHUVF
xBtcrAdLA0CAdlKU/2ZM/0nvMqKjZjM41vT9T/1CHgJ1EyAFSKP4L+0xt93FesW42Q2Tj2UA4D8G
OJ1h/IpEAv5ko/dpRb0g2+MdZvo9wi7xKdFCXc6lTjJqVAXEZitCAZwbZb6vmRu3xt7411LZlymd
wwKPA/QqaQagK4gSCVf5uUKk4y+Cas7VM7/BXFx30LmkpZzh2nq5kgwK43lEhT3NvTOn8w/WrvTU
j4XH5z3t42i8i/sHRey2ZGjCgkO2utluAjCXI3Iu6dA/I/OtS5PCFyRbsdwPgDnK5OpbTxk41y/z
ECnsIS2ztxoYGj5nSmTqCcQHusoHb2lc56fMN8u9Cj4lW7qfB4uuqjkuEqrotXPXI76vxi3Hsx9S
Nb9b0urG/WE/pwyWY8Bl0Jr0anscjx1DRI026GoGyYFd/XasJNeSoU1HmIaj7SVuERA5wBwJaJco
QOlk/FIV457yjnc+ZXmZGlFh+/f1QLyOnQrmGpHbZ0bau1fkdBpRnIe5+UUoy7tF//hut3gpMGdq
YhlcDq728RSuS6kilqWWUz9QCwuTRfgcaV7SFGcF4lAa9WhwZNJMnzZrFB6y/20GI7fBmnPNJNAE
yntVA/BPCa+TsLifSNTh20giwnaMlphCrK6AznjbAyr4DoQsLk7om4muzmvSzmixjeI2pn31a+73
0Li/hS9wE7cfdZ6PgSQR6QlNJjUzDdSJp3BWZKFdW5q1a7yodv2ThPKL80TzoL2a52DIT40O1G8R
+ZqZfrsUhIW0ov7OPJUqLEjTpBsgO337MtCQ9x1D/DvGt7YoZNfKCmvGz2uClNj/im8lVJBO6092
gMk0HEaBZMZ7mhuKU3OXoHGL7iTNKlpHqPNBUoEhv7TAg5GKNK8qha6AW/9BNtvSd2mkXAGsjwix
0OughUoYF/z+kLRihESBGnr9j8WisRgvN7ROziaw9NRe8s2uR1UhMf5pIBi1O2AKLBGn7kYCzzHV
Bz3xaJJSQEmijjG8TovRWt1DKEm4TBGh/PdWeAqcOZSSH2yfaT364bxwsU1MkwD1h/k4gD4JlXNL
y5u5T+5lWUQuyQlIoIxjlUW1xx+wk2yzjDP/OA/AC1c/7xrRyrqfmzZUu/L2CcdaoWuEpRdq4Use
gD43bQGg1SiDcg4v6Jjdl95defvWy4bgY3OC+QzGISGuXe2+ybfPglpPEyBfcujsCrC1A3HMZDqF
WR0QwT0NPzQ0P78wdwKgrAGN6QqQdjG3ZCtRNB8JxhhW4p2aiVZQ1oxUxuOZ7mVum6zEN7PwpkfT
buXkdRHK0d/yCWdGAxDsYugU8cQjbkaQlYW6yqaSQDkNmDJ3fgWT6GJvJliXk12gC1oIaSEjB0Ft
yac7q3qTjqRc2JEidTZsvaRzH1dK8obBUpiSgGOo1sPguNY1ZBVO3pMhO3V51ohXxnKhX/p2plpG
/t23BMej5czyya2kMWi60Ll1m4kAXYTeOOlF3A3Dn6O2rMPCE2p4XxYUrl1h4k7FK24Pg/pdxgeS
P1Ilg8vt/slTvTGILWBAkeWie1jKmGj9Q0TTOPJfajY7M/HPJQ8ckYHBdyhzmyyCLjV5x6K5SO5S
fQ93MvJDdfGbbizJ74kE3q2q471pOdqN46v8invPm28qxs9W7iUDQOkKbQjwMHdO5Jx8Y5WHPkAG
suT1mMyaDvkjpZoiI/e3cZMSSIkF39U867SWQXR9M9tsp74m8Lwxq7gC456Oc5R4r5b6pM0M8DS5
N26bCU3b1ktUELoFdwo7TYth9oZ8oZIZ7oZIjbJUIJ9IUy8jraKI+ZPckz+1jvFvBfPCyO5TlVlb
Znf1U3t3qEvDKJuWaKcmIaalIabrbrbITXvSoih7wPsx2S07pFNuR+2VIYBfpAhiJxzl7OYBfQ3I
MfWJfYK5UHZPYyAdj3K+w0LF3BLNl1v8Vr9JSw/XY559KFQzp4TeAOuVi1hVJhmI6Nw5Eg3RycV4
fK8qpXDlp16F7wym8xjdBvYuPIDzKFfOxrA/mTXHcdNp2T7H0ukgOPqGZFSFxLZcTL+VVItZD/BU
qpJrRTdCC2Cgvg7c4JceBBVJohkJHpdBQ746MiUNJOijURMTyE8bCF1ARK9v9VAgIfNtZjgnOjuX
l8fA4wfqZH85yB5ldVAbWSTcJ2wUC6U/6foU8/X9T3U0LcEK5dmMec+Xu9QBeggzKswDfY0dWlBk
XHoI5PLGIYyPkn3DmboIZLNaS4cLbAt4u+b62b0aURDIzRUy1FNa8DK5V5W6gwEswq3576iw3Qwk
pK9PhLNlwB1FqXSlg1ntuyqGWYQsBnz1o5UCQZlkWGlKc3Veb3hv4jK1oYSH7/5ZcVGAINj+ROCw
nEzCUf51seW2LTFbkDk8Lfa5nyEwwyJLNAWnwVxjeydPBJudTD4hQ7KmC/RJUIrF+EW6iH4eckzA
Gyg+Oa6oUd6fRzZlb99tHbJmpjSAv+gZXDNtYkyoqOIlDEBr/ATXs6qqGDVmH6OYXBwiTsPDCBe8
xUuRi88HbQclgr/UqyDv+sUGvJXmUyB4tIZw4hs963WnH7LvG2Dfmf0s5kwBmM4u7uRIg/rXAMrk
9GzREKXytj8xeKxkw9PMXc86kbqvvvjS8P6zV/Drnvi+NMnSojfEe0waQnaMaUCR6Pt05aYv6DxK
wWX+t15ND7AXU7G0joX3GnRJEZ2Ehxg+FY/0x380GnC8GVceZNP/+M60Mz0vb1S92GVE3ZOEBeKq
/6aPKYQtDUPKh7EEOP74BbWU090eoGuebqVkUXq+lJc0sypcIBteuaTaWK9Js68zJal7OOZslf9I
8vBIk96fu4WrUmziV+NIQFeFGivoz8Djo8f9+LBEzMZgfEeV7QKBBI/Bcm1GhOhDTBKRWNunBlwB
bl1n6YXD1Yj/n/ZCXNG21U/t7Rww039FXkr7GNrZvPcz3QhK7mT2M2WBfFO/9osj24ODIIsNWnoe
daG29yPGkr8RdJpRiLFNE7KW3Zvo0fbe7JxrtdXv3aXoNMWg/TyrAVhf8EYGOwHF25fsFJg4Hh55
+zcfS5K42Hw5WJ6boDMiJfl6cxx4uiQ1DPilr9R/KiNbY+uAoKjW/cVLL4B7R5L3G1edD/o2iev2
LVok+znsYaiLJCBQQ8WvHg3Er3LEJ+c2DB5EJwOvqgBTejh2MPbKia50kffGwKpsq8JKMI969ii0
/qJC8nnf/svqI7YOrkn2hwLj8ZuDUcrkTjiSRGB29iMjhCtGv41m8Fiwm04bMVU1BQxwHyFfhFPM
1qvRrJ4PSGmJiqNkwtvoxxoH4Pz8B+Xi9/3LR13++kRmBpoIS6K+I/qQKrOh1yLeW8BRYCsqRloP
bBhQ8vsZbJjYcQ5sx7+/GjEMxlwmQZ8JAfIjInTphfFUFVgAib4yUhBryxKuxNjFrF/jNe/MesTg
LMh6nm3fwCSsW1CHbIJuNeUsV5zCHQmhSPOr+TQoOLDF/KB97jOXsU/mPK6UyL9Z78u9p0mlD2Y2
niJek+XOLSnWd1U9mg4GLybRkOxOeM4uDckxxePbdNBJC/0gqGmG7uPClL5qPI0MD/b5FKvxvv4/
iL+fkca2+7DbVen1u+7HGfAsaNPOArmlDSmCUNhibDfTPPTAhdye4X1rdaVokVXMvu4ztJMWIUd2
EWVFiAT0LvjkQs0R93da/T36yn63QocqvitoDGB4a46XHkTcOMidLa5LL3bxaP2Y8kHISx1y/xXK
6vA2tnyvA5FzBBUC9/fO6bVH9w1OfbSMat6Xrz9klawdyA1QF6VBLc6bDC55SlVPUybIQEQ4NrWq
nb0qQxLSmugBr/Pk4HCXS81fFLzxTBUiZRai9rJNpxPjXMyiKz4FKyYV++QOeWCpEzUD7Mwor0LH
gSlLW6BWvLGaIFjv//Hax5cx0eeePyPJnCpW5SNHDRTpDigihebiHAmYMhKDZkLuIlllPTktvqLp
3PdUJosr3NBzGTDg+Rh71GKHYWeqJsuMRxTfelX+Kp68vsC0pHCk+As0zTzX0at7TnoqVAs9p68/
kIa3mYE3YZlyWWoXojKvfPCtCDD5KqyIwpwv5UmYI1NyI8cRWmHv26S/bMMmRSWGfuwxulsRN2ao
GoaCMF8hUwVurqe5DmQ5EQNrY7opwkyfWL83WQMie3TgKLMp4Q8qMrpHEmhhC13nstoZAUzQtobm
IY329Lip4TQ0pm9X0L++V0taeuTV4DBiwxSJSLO3hoGoe+uxMOuZStqg+gmSNfTbuUm3WsKhJKWz
MWWn72hpQWN9gG14cCbZOg7/OEy5AKIjZb2BEDUGlraaeoxQPA/fmAZjDmw6aKk1GwIMj3Kj3ZOx
grEfCasTzvbtWu4W2KvA+IcjafgxjkmH0tGLJSIm+W9KkI/PtetqZ7bHxA66xi29NzB1V634EGa/
6BsuWZrjIpAKCkv55UddQlSgvgYRWz8XFJpCmnpYdvTKtpBkdjJ4+OlfNMYxnr9PFknd4KahcHSZ
fcyp0heKQY2zbhfFx0hIBDp+Dgep7zfokjtPAurN4ti2RiL8SHL4YpRitBcA0bxZJHrochJMTP+H
DsD0ckHrJnLV/3wxVfNieNCFElw9j3iR7Sg58MU1SQcMOJmoYgyIUlpv/CTbMivQfeD5EKuYrnka
YfPaEzfaMAQuG2dDHtYij/AqnDRga087fsOp4xVzsB+LF/M8nVjaRLuY25wOThtUh+H6oDShJSnD
AxW6Ug5vNMRL6+gHfz5OuYYyphlwxjfDF5cplo+pdnU5kzi9oMPxOhAwnr1CJZIBQL3OPtIkGivW
gZ8WjJI715Ntgo9n4jngDBZ9Mprp7rpTPvIVeo5pL2otpyie374IjJiewzEAoz0eRUDg8HhLQK/x
MI3Grg2ANnNIDOVkzC8RtBquB7B6XRaC7yU3xN4ClEF/NdKeZZoJh52QAe2U1RU4mgYh6GHGTKzX
/9s0JJA4WpPqAtOlZh4VQJ+tGigGVNM8KPKmDOBxZPlJbiW1VJwaP+exi2yISzCs3hMocR8XbHTH
3+pnRYoQOHEoqsCy4dDus7sMHS9kC8yto5nMjhkDXikRTePMia0cbZSZBn+FjlAjpCAUNRpoZCWj
Z9naCiKN3hK6yckz3AgBfZijWPtDkKulRWmnpY/+92mBgaTQnVgjpg54RGRZilq1KI4gFCD42bRo
hrEQrVPiZ9DGqD2zivJv+QSrs3MJKMPuoGTZNZXUprHDCU3laDJ5exNrs6Y4oiIwsgD3ziHqQORW
MnUTwLcqO1PcMuAEWrRUhKYtnLJQSgqw3uO3rrwsQdoHRiZJUqjPWqv0yX4w/OF4fDwPrrMuPlzl
KHhn9T4N0OYJ92C4gAQvED6cx5l2UP/FzhQN9GP6MdCFgoeLCUPDnthoGLvYyh2xQOaVAgQd+U9y
mclG6Hahn4dOBS/d2TdGEBkFhhui0h/D7qizJiuS3gg2b82DAw6Azux40L7fqddPm9K+oPWO6V+C
+Annj9NGYchlTenHjoOJzLSaRZtDTM2e27EvfoAsmDeGJGC1HP9I6vj5V7/5510UWYHEtQk5ihUL
Z+01lLWs+JLF7DjiKnYd+D3pOSVWBlWOFoNa42N5HYDfRFxdkvVkisLYdEZ9QJO3QP6DwV2ZiKI0
LGi1Su/pfbPW982MV4Irhzedma0BDc4LxOrbhVvcznk8KzL15GQnAy8Efel1ob3v/QsinNS2A9ae
v+TLw60/w4xxrd8WoRV3AxHaMPz1KwKu0+r8+F0pYndxg/d4votwN368VS4wawZbkhejRJoM/hh2
cPoAcszZxcErP+8L+q4T2Bw56VWmbispmydhdghtAaAZ4gvRX0qM/nPH1rBYh8PJrl0PHUXcdeNp
FRyF2fcpovLy4bg0WvWbbvieu/0OE8Hxz96Sbm8mL50CMXxcbdXz3BCdQn27+MUdshwWu9qBcuC+
npj6tyorSS76HB0N8gFfxTJerA5ta4IY6mTAO88TXPKZTLrBO3fCIlRSNfC5pQmEJhTQ/RNn+n4r
AH2s5e3dtHL3uov/X8b6piO+ywEnytSUs3gKpp1o+QxizmRxZHmhBhfqxMziQQNhDVrqhhIt9Jor
AOzSEFMFtGyTSrOpXgkuy0KJsK3eWWcHYxRNEfQCBHbWy8KkmkTpWJoemCPsvB/uUp5ZDhNj9o68
eMYqS8pwrPLv8KbxB47UPVxeLP7spFdQODR0vD2DzIvm3v/ox+DnAbbSl629TE9oBgTwanmWMUWM
5EKB4UUigRsX1uFdS9AOPEi23po8dThiMWzvh8gOEs47qWHpSPGc7WUxQxWURGxBxqxtIuU8AdUh
+0NfuOlNhNfP/Ld/h20WdRfqSB0NiYRGnVCRTXsW0JLYyoTRHTuJdLt5N1owcFYfMeHqAEH7+3G1
GyAZwlMIvoLmW6KzWPmSqT07wRJGO8uvgSP2IEW9yRw+ZmkMkP5lFjreaGcnSnr6Ro7Nrpx+HccR
V44m4nunaBoNRwyrc/IUAy893Utwiov7Y74y8p1LYcUuLqb8b4s2X+mQp/mpw9xj1w7vWknTaWEp
NkuJAqSBMSF9QsaqufgGJGqZylSAxQk0Id9YON7jebKIeBfYBDe/Um1IbnvRgCvIjNhZvnXkOx3k
HYYoZOYo2qxLaLzfHy+pMVohuI4MZaHeVof5KH6H0T8mLnjjK3IgY8qjj5T3sZoMk8RmJuHiCT3M
tfeHt49Fr6Z4Kegw+tbEqZ8CSPUfO5Up/d90SEyiR+dh4kzvpU+nHD5yzujoTi9RNOHFGR7lSMd5
iLYf0yrM9NnSnf7TSRXqXS8k+dpFg33ltUNotPkwI8GwuKcnJ+yVQahrHtpkvIRWeLPP92pYOVMj
mIS4gxPyeK1FNO19DVA98flmzqFo2z4B5+8r38ld7jszGX7eLMyLrg4Klo5JTIFP1XxgMZr4TwSC
e7JvmGqUK1YO+pgCAl/6bz2VWrRZSqTPm0InN4a761er7wu3YKeOvhFLmHUQ/hjJYYqrotS0nme6
y8fnpy1d/7R8MVp0FzR48BMJ2c/gZrqd2rvbsOJPClp1/PiztsOEeea0NZxhedjC6Iu5eJGDyXLQ
y9lmUh1TfrcYLxO7+tP/NG7u7mVsT/Xpqx7PP1F/U8M4Cgxoq3hK+dqn+HbS6o4IqG0m7J1QPCxg
EZOCWkfuXhAcBu7ewNVu4cjMxgqrMU3Dl2EFrLBGQv2dFKMTuM4ltjiZh9VMUxTOZHauyrh8mLz2
0AeXahrc9oSKYttOuBQWnVunRRWZlh4NXIO5A7TWFQgRRjSe+9qSgw1L3z8TyueazKAaSMeUKJyd
rIwxMl4ggKmMEgDDlNSsjoV5B2/5uAcFvRas3FdNS00UGRA/NgWz1gj1DrPpDqdLWnpCxxMK8iqs
KK0x/3ID2QV7G7+nL65VoXcEjn51gXpix0AyKp3n2KS7duvQnWNDIa3rHyMWVE96oPnV8cBbqBXo
d9d7IFtFwQ+xOvp4HmnNeE+8MpaZmLLgv+cVe2mlNeGGbpXC2kWkf/lJfWHJYUy0+Nlwif89TIts
eudpimW0vBNl6qU/O0hLdhvoV8RjK+x80fVcOA3VAjqgszCrCrdBaEd6eL2S1jtA/lB095XjiMEF
zoGv3zdFkJkNIH4lt0wqByn/WnkA8TJ5C1yuhhbZCcZqC9YSNSBhqJ2+2+CkSnYIiMhP19m3fNJd
9H6ArYTIAtGGfgiDK/AM4ITGoETn76SACTQ+wS/zT4NLpptURXHNVFrKVEiYvLs6JppavyW26APH
NCPY4cZBLNRfxR78YZz0C39MhwBkUol2tvJHEwPTqlPv3pq8mTG4StIA6/6LqLdi1/Y+hXAZZSpN
8H2bBL1zEmsZN5lxTy+LrGmo/59ojpO7u+LpSR2WH9jhWmLOFHx9fhYbIhF0IY1HTQVoeZfF2DAZ
mhxRNLpDUD4WTUy4Y4bOXnMj9EAYwySKGj+LytzFeQHR8jKrouxG6QnNWaBSnhnaiSQ8ca4OP4L0
pM4Qd2Bxpfagp59jGxh0V9aUW+j56u+aUlFJlqTPUfxnH8oX+/uqUeTnETCGw6hOZgm722hACGg6
WvrEQlFzoG7T9h09/sYNg6n2+Lc1u9HWKnb4jzgyKc1becBcsZJOIPwsLvHHX0cJ5dLQtO8qfXrg
GX8uskIlGNIbJxMs49tT3nbEGNbXsSbrHz5oKebIg+UDmHKxm0W94D3nCFtOMtfbTlNEBWD+4wMY
lKElHMnzFl2GWpbh1dHS8+QRTd6Ughn/AxxoxLAykpfKVOdG0JrVBlGZoq1hYHvD0vbCda3noQlK
WigqA0u/gPByIAcNDMVH1OIcSaEEFM6GcEsxAY07W2inIcE0IjmfzQRrHyLKUCSUtEZxzW8BeHeY
ddJMS+p/HcYO/S7LpsKAAAzyatQnLzMVMsGXMsCcBZZobs9VeoqCd8GHnpQ2E9DyWsN85kvvIlBd
HyF7BKVYoOF2zIG8RYYKi1j2Sq13yejEzNqb/kKwufqTtdLmq0tqECf1O0T/Q2lJbAqFYmUqtror
q5+QveizHX/Etoi2x57nS/KXMLtfZEbi6Lzyd5q2/UXsLq+gLCX5C0C4Zm+vOy4lfVuk1oGBQtq3
ECRGdCmcS6TREKnUyJ9OBvNCrl9WdsDbuY5jJYnKmqVcMem/QY3OAlPcVSZZAXpefIN+U4343izW
4wk6qLDN59p7UJQD857jhyLvzbMVK2AKKeAsduO/5P9nP5dQRGk4p87XlAFHIH6C86A1plSeVuh5
OaBBrnjHqerIJUJ/BNONHewUBexh83VuTKPJCRx5QpzWIabh+Og6hxFIGEMvNeCWi2Lgm0sFnHMV
N4qD26vnKuQ8zEMlNR4XA0iStUjRyJL63ppnwUGHx0pSO/aPaFMatc81fpl4E3hexCo2dYqCyMAM
oA7Lhvq97P1goAngkFcmGrRlOu2ebzmZoMMYGr9U9okv3D39+55xdiuXKlWP3l+6BsVfRfQytpg0
o/fD9V5NCNcdyBb7ieEyVfKUxrlZjMTdU/ANA06G+volbvkvXGsGC9wX4ysiggkcqSslv/hWD+Kv
dHbRyoHSOXgiz+5NYzOPQ6aNX+dl2dkBgzi6uWcDwzzMPOhfzpZP4zsyp4qFjyaNX1XOp93rcz6E
j+AZpg1QKBWjHyOQt/078p3cklcdS6fk9O8xS5ghAXCrTNq15VP9Ym2zAPej6+cwXmf3qP3I258m
Cd0Sy6xxQNlFyLsixMWukJlPf3zuoB+G+lYd1PC+aBLj1DHyhWbIt1GBNhOdPa1jXPLoodDJ3Sj1
3d2mOhRT+aU08imDuyx1gXwqf1AkbN9sjLwsmQGkY9XOknulWtMscIrsEVvHnRy986GysfCT2JI5
p24dru0ZaM+WKTm/w9Ygp3gfIXnuIYB6MjEAJ6rB3//XPBhMqIftFnVCFMZxqgm72FaFjEMAmSlJ
gNMcOj+R4PjPduKG4K6XVbocI13PN2Xn/hdC6ZzlA2JqvEbsCAdM3BpkoXUGL9sD7fCgarD2xnUg
vHL/1Gsa0JMaD5/pREsEmlq9M6xQ+S6EO3zpH3pm/TysJKpMQGZbzTgWjPL03eAH0oHPzbPT4ZPL
h4Y4hFLlwoBOZDZ9HmKu4uP5nIovBDO7ETTJv9gArFr4C6c94f3HMn5vsBWlVMicICRa6Ee/fqdk
0VUVv+GmIIIaoNPOsW9VUHIGAoG21XyzskUuBc/K6n77Fbqc7EL5Lei/tKXvtsa4S8G4/rZdtkzm
FBAjPD2MsBtZcQX39ZiHXV8qUWGgk7d6vinQ8Tf58FBqGxEjaLgXTdigy7UEa6IhXegEdh9/NBRA
ELXdGWZSsc6QO6rmttgf15t8bDBza2+c09npTK/lVXjNEQzXFCZBW0SdktSmjrHWtPM2iNrw9xAB
iUFmiccsQjewrxlYY9trOEs058iVIEma0wUo1lf89g0b+V1R8Ew535yusWT6KretLBfoeU7qPmGJ
SSpwTvAe+RKrO20+rnz0i3jh6+8M6SGbbCSehZOt8P9aFM6kbpImGPOT7tyt7EOFTmIpDMNQQGn9
P0dw+H29mwBNgRZ3gGD6p80cpDaL0Fcvq8pCVo+QP0iToa3oqllmoIV2ilrPdESweVCabgsgJV8i
r8NECCsVMmh4ECt0rzJyTYAk2YhvaXMosd8Za5zDkKQOV5Gjz0CDcnKqcW0dLeQX4mPw3ptx/3Zl
VHp+lTOi85YnEdICDdXWyMMmBkDhXttgrxf99Sp6nz99gZjQPDyiTmQR+g2ZUqVhioTQPAz11ad/
HMUCFulWgw5yAOVibn2N8yNghkH4LRdFZpHLHcnw6vgdj2E5bkVMDpU1lXj2jLo3EmfpA4dMwqWC
VPQO7cJ8jYjibbgOlmgbTF4cKNKBysdRlvod3DmeTSyVeeA4KDe/vHPWJHuOAyOUTg0yUl3OBsJb
RuuZlkPou7Lq7V5UysI8aYY6ar4VSzuuQM6+hCfUXlftWRxAB1Z6+zplsb/ydLr4CJrliNnWBdNH
7XUfVIPZIAt/GVOtZRDEeWk715usevKHYcEKC499bUCaI3X9C6bR4eDoR4fKZEkTvzjpZ9Zr45OA
+XBvnOzCEKLc956mX5YcIJMV49yyRJNh9syAdINTcDSbTOlBWy7XnvI3KZrhCusvzJNcUbHAZu/M
ifIqgx4d9YLtaTsmzlF3xOaKYA4i9jcReKMTzVYEAZIz1guLdt6v8LFv4wVCgAHXidp/4FHhm41N
EuQrzewRZ2sqIjShcxcUV3d545hEuXNM/PIKGghXmK/WEs0EX/HIMPs2m3ipsCpGut2Vlj2HQ/n0
6RGNNBmDdzpGakx33rno0zttKE/gagVHM4I+yzYVrR4AqmZ33+E4aMIe/4RU1XPa4RZQKeUoXfSS
zKpJ+sk2XerI/VyGWWMbAMhX2rQmsYY0mQvFwCvuCAXtK809fD2PlW1sGoRmLIUG+aik+SVuUIB3
rOum2TCDga/j9+sw/AcuIqTyeo0x352sg+LOkovC2SBDZJwXBYHA/LaivBUKw2tImuZyUZsCnG8K
9d+/7MwFgbecAytRmmtqLQrUXdR0FiQ7t9weVzY/M1njL2SEXPHsWS8Cjlub025KWanQqrE75k8y
+NWn1CxgGTcSxnKOZr/W3LW90AhJYSZrqeaHhtUOUAEa0wSVXKRZJJV9AbfLJnvWCmM645ei2Ke1
1LDv/rpjx/S4AUJkNmDFj5k/ljbwk+UKn/Sp/H0i8JMgnWjPbWwF6QpvSUG2WB2x0HS63yjnVw/t
wfO7h0OZS/L2fWcFw6ZqogMpexwLPq5FtD6mPUh6FKJT6dj2KIPuDrb4aypRxyGSoGGF5NQJAGAS
h+4rppwxqo9IuraTcBKRVC8wNfuS6fSeKLc2oOXE4cMtU6pUgfnZvk3XMsMINsaedPWpDgoz+WDJ
r0t4qtM3K3TzEwuLLeJuBBlO4+64MMjry5/DO9CCbz4JOSO4iBq8tK8x9X3pro42SBYomwE6dQjP
hLRi2E/FJ7jo6LiJtXVdsZW/lY+Rbpjq6c3T0f9spkjgHlT0GCMqgrR9GWMsZcC73j8DyGIFTAVp
ZXu7TREc15XVOYF/OrYOHLrZBUCM7DzQ+9SvZ1HZIs5x/oCJJA7mN1BJ1ShMLPrxObISXdxQZReH
jAHah85K/VwCVE+IJLnzvnIxaF+O71eK9TBKDBNS8zgF3U89eMREoxTZyOvKB5Kaj62in2BZ/hqQ
YKC3kmWw7xuoMkwjn4eGOMBMezNstVvVMTz+E70mBlBACjg0LPVEewKM92LfX1B3YVZxqU7X36mz
oCqsHao+5gpO6P1i675hqaCnYtuoD3481P/jDNtVHd91ck26Ve7PBOUKH7Xk61YxhEis92oDAx8U
M0rSg+RVs6WFqPsrzETWb+YEp1deBp+dYuGp392LvfQK3jZhg01yUsXDhOv1HADRhR5wWZdCOfUF
14HnLx7t/zYn+hp5rCJjaLRSqXr2K7kX9QDR2VSnhH4XvjLDC9JCUNIQeRvR5ezYarwlUsa7/jA8
wy2MTnLEQMsI+S8voazaNYo6CgVmRwguj96OccTMt3MW+Eyks1yQnu9j7ZnxJqPRhYdr0blBUF7f
shTfSHvfTIdP6Zm9XctCucVFF+NtQjLol+AaOECjpEz65FrNVavsdZnXJEw91xgOqWOY0qth41Xn
HgNuy1/AARr2dnuooS/XeoHLO/AKsgvBeCxLGINSHNLqvW+04xhVB4bU/lWU0K08ykWYMzpVCubY
zIuzsUVWD4zT6kWJqmX1gpGk4xAmNuMzSachmxrjslvN+deIkBy50+NK8xyJJCtnfEWCFgs3xOHD
VeDnX26GarYxhtSWI7E5MBjalAamFpLJtWKdDZ+ErmnIjg/NG24RZ9f4Koj5NGVjIgB48A+9hyFO
pBBZ/ehvzWEi2ctO4d7GZLCt/cDEyKnZZwZW3KDk/Fy9upBDnVRd6xLKcWKroP0J8VfwSQ7b7gRW
bQ4HaIvj/n3roVGPjmA4gv7YqaG9gEGBr2QtTTWfogB2BTD96hYc0FPrPyTRyqB78ABE8YmRiVkn
WhG9+f4ARX5VlfD2UEHkJjnUK+y+ofj6diJimVQoHKmRu5Kiz0pWmkp9AMhKCsPMmYCqiZtfhpW+
LzjIyfoGcAL/wWxxa8NEemDtQvFgo237L61wDtF0RGvOj+Cw4X5fIhfgihj3VMNuTETF3WQ+FVzC
cGAOMlJjnadKTxz7iioODvPOn+QKYy3qYyphwRHCXOLaQWJoGmxrJWicPbeSchTWNr/TYV8Iwr5N
3gaRhTubjDCNgK3Fl7GJELhuIS9/KMysqOi9A40Tgyeg84UOoJVwJYK9TPCXc/0THwdg63WSbhKp
NqiqTQBXp1vuABxIMthAmPYr7TVQRJvkxZROFSRzMtp+H/YfeuCz68wl3vflylidWNw8ngNtiZVl
WfAoSvdUDU9flyevQ/+IJWg0hQTiF3NCOM1cmOORwNAazGrdB81vn4hRRH34ie2Beml3xge+XuJ7
9gasneaLk4YeMDHW4kc0toiUxfP3R3Mk41ZJ1v7Q6CaAHEeyDISDJ/lQdOUbmpHfTmZKujo1MrR0
zjA9CCX+Vzwdx/dmXyGnpCYbJdTkyuKZMdReBpQL2xhk1DbEQXpjRhszAr96yWMyjfdqIOi4xQUZ
LddUEgf9UM3hi3AC5juGMa+hIIq3W7dKxwsBoRvn59ln+IP8oh49VI9//9Ij8xla79c8kRXX75Mr
MYFbokqwMe3ZQGx1nZgLhQ64X2LlR5s+rbZN9FdkZQOrWdEUjBi7B15bH6+AQ3bRNV6rvk0DlemO
xwNoj4h9yK6tLOY0RVFP3YePlloVhIoCxuolU1ilp9pvUglwt7+n+opLEQUxMh1RhERUilSsYNo4
oJ2xSgqJkB5O5sSRg4LVHhTf30gYgDE/ANJtsljY8tP22yVCS/MMdAOA7WhQPRbr6cVpLNJsKOo8
9+wjK/OrPiMhIJEsl+VgteU8m8vfWksEnnL4VxilBNrHkV8ChOgURy5vlplTFITdLHQIeGmWedH0
HXo7/l9WqD1oSL7Kf4bp9FY/ci5dG398BXEIf4q/o8dfphoEEa5MRq/BSFwV/bb/0ZXNEas7emRk
x1BzzEk4GlybodwxbyTrAQNK53jwirey2JPqrDHrk/Dqc5yTi4oUevjtwJD7+gQ5+rVW5UkIGpJ2
1jJqTMBO0r4x9Fa9SeegPXafD4MN8sR7TfsH/ut7D2cnGcg/DxMaxSm6k6cIshBbmaw6v3MWqkz1
/+0hm6TIC5ysM35KLsO8kaKkLQVi+hCSfN0+DZayUW5tQHpFWYrfS5pPcK7Z/wmbr+XV0MhjsNu+
WK1x7KmUENX6FJnWTIOhqtzq8KG05wfMcfOWq+RtvLbiC8ycEPEJCh5fxV+Di+5q78tHUBJrtBXv
RS6kSqjsmBazeKs2vAl2zxTS8ISSkTSwzuybW2EYuFTGBSKQ4SBck1NSt29Nxi9nLDqR6dmD2AkM
ooYFzKiyHRgAY/efE+x+oGoAZh/NhAJ+3ugKo5BOkXoAOjjxS3MqlMf2A0zAZnkiG02g3sxztDyh
pqrOt6eLG2jnjoyqxbLJdSS3+gqIzVOSXlrHoq68GHmknDpJm1LcpoRjPSzyj9cGYiVla9tXyY/1
Q/E6xcOT6oQ0t55psTYgQrRULUGN9cVYw/Ez0bDywBciVt2yKrkGw7r1DXxQ9VwXyG/Ylj4Arz/t
xboMDuq1GuIpOrsXxiyYKs8T5cYQXkGRmAKWjBO2eGyF9BN3uGKm0lxg7mA4TGZIvUL9FNwgcoAC
FXNKpzNonrZrS/VGpsMG7wmYwFyRr23jPq1L7TYRnnO2sp8Wm+iCIUktgFBT/VHc4NOdX46GRHjm
w+3ZtT2bvHjMC4RB9kERhzDjimD86TUkLG7EFoqXR7JsTvwB/L3eHEBxjfwpMifcR6VU8HZZNAgR
Q8gAVKJOOYb/iac56/jLtmGVNxoWsnusob/YSy60tvj0okXMt65K/Q3yYy9CARLMF8gE0BwfVHIn
OHb822oZGB6jWqv/yw/ssbko+hUeDDBAR7UWAF2Uin0um2xQCLiHxue52/Q6lU6VSn37eBj1XKcg
73Gp2XZXDDgbkQ7SpPSfiwxHEqauo1zSytgaSrl49m618ZuQCsWrEYsT3wsQ8MBeetTgd5+qc7tq
RW0qkyf2y6Kz46UTLwx6kattkCXj51yoo0UWWvNvryJV0jz/KcK29VMF09Rz6uj14TedKfzZa3Zj
4R/QwmIRxJQTimjZgp+VEhtXWhW1zzhA+eXF2479hwuML9Yt7pBb11moT/O0isAKzXdOl7xmbMO/
teRzOgdQRLzYcP7gM1rKRC7csGt37dAVO1kmQ0lljbiEXpiDgEh2kCUhoA4ve5rPZRZjarQ06YrN
RO3hlWSg6sfGPMRN1Ite7VmdOzOcDdQcdlFDJltch/BR4kg2Dhr3+9E8VtvEp2f5Jc9VCRRtP/i4
3CpAandxQ+lVLmIVBrr8LI2w5oAfdGNzqbG2ISa/vyoQiXLYI4nm7Rhh7xN7dLvz+C/9J/AYx7Tp
WFsJWDsN/M6BXWVyx2FxcWH7E+bVbkaQOXrH36dznp3OC3X9BSq5er/T6w9qqX8YJDW/2V+5d5Mk
wBkGqaHA9kLjEcLUuOU0sp/x4qYB8BOJ0PuVTFOyBsqm7+7nkPXHf+Ygm52KpO5W90sv/dHQH7FH
JNJIQGz4HMAJ3cY9G8dB6uEPJFL5WLRfKueXwzEoI44d3OszxRa6oEqf+xWvZupTNtnTtrnSM8TY
AfQHOQHFh2421XzFYMvdWCAU1QK7h6/LXAz3QjBrQOhxWxairLitg44iDvWKdXLqCzvITVWv+Nwc
jPUMcuR5OtlPL/AJLHS7FoQO5nyDrdr6oWtwJddICTbNLUajjCzljZxhk514MGAkIIIH34IzEKIO
EJxCn+/p/8WvJE38cGIc4DAd5keuLBCTdpEG+7UpQsfD2sFu4OUAovKjQ8hA0rFDlDNHDTsyfQa4
h+vJ7J0kZH8jsidtbSTZdWMh5rPLUJm5CpLO67qm6XjIPH7N0f+wteS84v1awBvsRNc4e32runmh
xy1lxLIcU6/8KQo8rSbFNtm/NkCZajCqJS4Iwr497saYPF2rQGS2BmKa6HWjw+k4Sz+AGRm95sdW
690ltUWNYA06dJJLk+TRjQDJ/iuNJHGQgWKChlIA9CYx1h+WnBDCTuUNw46crtdl20jgHAnCD9f2
nWTZuv4HvidZW8EgYFzdpXz2Q2f6NZEpRXFpmfN1tBrKyoRLxJCTArKX3hIeWCywz43GFBnWlrb9
ssOc4GhRn4vNhvxEl0IwSINl+Jzlg642ium9Wf+AA86RAkaCWHRJHjj+pbrdza0oNQ8z/941tYrU
Vv/Af68J1GXEz9TFw0xxH0pLsolopallv8Hb3WoLV4bRwgqWB+jNFHOG2l5DYExplT7ug049QH7P
hE7jsAyDSML7seQCX+G0SFftCQy/8Vqy8S+rnUdXUeIyKubnmWwSNrqJfgtXu1LGgsRWmuVuOe/6
WNtw8spxWfCtA2HbqayE3x1lRy3Z5XJDHY8FojXOgnqTMir4KZilCwdYU+sauN2r9fq2nd0ypFxk
GHPGqe9krOzsDjuRjdlqkEKCBRj44g+PJ/7AUH1x50jsp8V+96viPEmDFBqn8eyjhg6mW55lCWuP
ryDkRPikoAH7RfyqAF/Fd64TREx9no3RoGfLqQjC2rpCyY21RTVcfviE8/mwFwBrCxB6qEtbUkje
7kxXfKQPKL/T6IFv/mJAr2jgux+RDxD4/miCvwXNmHl9bPhR36zfYtYo90VXePjykS8XYTuOb2fn
MMPdzvFd8SiBc9/zSLrNxwdy37p9sOxdSBACHdtE7v4E1+a+phSLzcq+TJ4lyVmeO2jyVxcYxAxr
IKGqS2wximsrryPvqFPTlhkG4sWR185skX3GhxsrjIfbDxtgZ3WxNwKpSYK+6/oA1Nw6kr20ldin
IMBIb1V+kyEXrYaZQp+cokx+RI+SKgbZKkD75jfVylsQok+CQwnigqTaAGkcoPEWHIE1WSaRTXFF
SF9jpfRZyRLpG0+0gG9ZBbzW2jh6E3OJr4q5J+OyltjyG5QXuAEYpjNSH8Ia1wERTArfble917AQ
guMjLqZ4Gn0TB8KKofyp5/YW2VBW12BH5ZP554cRVr/TpYwrOvmjP3vWKRTxYsB1an7+JKrmjfgX
WKYq/++VRBqnFtdSKs4NSxatrCax1Pl3LTDU6nHSQgKhanSrUK1rV0d8m1CBDvlfvMolCuc02gV2
KjnjeUB1cdOICc//Q6VPgeSG5SilVPklJ9M0HRNvclTpbLZTUO+0K8eDdgk0Z77bhiYccn/azobG
RnxIXEbCmRCzqFeu3hJ2gOokXomRwq03LIkMiUIM/oMqfYACnY7PrqA+rPH9xKfdCHeKtFd0zJIi
1q4TmCeDxCjwzQYdiISKPdIpYGnx/qvDcXVfMLSyLq6Wi2JiDa4teiELnQEvLAIMvSFNE9F4Ra/S
ioL9SIGA/dXceS0JXyqovl2TIebe8hjLgdv40WCyA5UlWkKnh4idOIl/fD22Q7eD4O/DHJDkrgit
aPBLD9CDGgTSDEnTfjyol8BrWnVycIxqtNfWekD/F4XymM5z9mCoDRV5CfCc31SprfStUPxp5OZT
IDzZKKYsRKPDYXKjlNILAICI08GG50LEYuwLhWxRlUjJ8kFnoH+gUt/5EsY7BgMMVGjjacwbyGtn
FNq+VFr2eoBejcnI67Z+SBC0AUtVtkB0oA9WW2p77o9Q+/RZ/qraUC9S8cwKAOeoXpO5rzmXiBqX
vBuron0i65PO2JTcE5O8B+ovt3iC5VBuImSYW4+plcwitPYHx/SImjm/jagKcNYVnFmvpq1ij+x5
4G+YP7pVUbK1y0oxLl1jvBuBhVk8K1FX9VtXLpEJylM/5WSDu4/VXNDW6GHzu5eCpD18kHhl1J2F
MbyAIIOH4FYZwuep145m3m/hJpA2Yz0ZREpiKOAAYg0vV/XJqcV6tNX+3o3whZCe7a/PmLng1X//
rJSLAX2DMdFNxfBFxiPYcjSsHknv3xYIMaA7I7EIsFVFhkcBo1qJZ6tP5H220h54zAU4JYNKZNIO
o0Gzv8GO6H6Z0YIypv4TX4hYx2WQ0bfoAwhvpkNLI78tl+yF/orFzobA1oYqcoSK9MACmM79GiLw
YUIVmnmoB7cqCFt+Hl/AIAR+R7S6L+HxqqUqXLo+sV1sX2U5gmgAWA3h3tzLLM5b+MlumBC1ONaS
qGzjylwcVLeGGYzRfZnv65WoJJr9c64Ailj0Ov0hPx5v+VieVaJp58WjV1jMmWjbKHl7e7599qLd
oWabqfydh6BLsXn4KBwdkfCbGAVChzc+1pqByhavvES0XJ2eyYlYTYUKF8itFwSPHdVFpOzuZmU7
w7c/NfP+suvn+ei/oDdpl/NPrY4hAJlXVjGFISp8crfzC0cevKML9vjcHMxy5APPuyKkBFoFyOfA
jJWLlrjPQVJhm+gYiGwIC6LADGtEM2gxApPSTcr4HyAnsqcNeq4Dp7PpvRDYxkeRdGSe5Z5Eavkf
ZlmrqWclLTfooNzPHBmi7duTBcniRm8cfF2pOoC3G6p5hbO4JHDhU1/BSm819fW8MEDr48R34MfO
CVBV9znqC8PsNaopp2r7SR7NQQYIle6YL5rUhe00Vk2nlMiiIArkJvsdOjSf24vzLVvRX3dw+J0U
WHTrJrWJdZYv1r9ythFsWj5Zur1WN9hHUHFnEyF2E0cthAx53eSvV0fkIaEaYZT6B5vr1YEBdFQm
0v4Abfp9Xw2V9jJiIotiUtD+nfR/rpsUsFvIRcqR/hNUdAt1/DHVTHuo3U0MUCwQKTfPA6PJgBEh
K/6FZCyIqiCNI5R2KxB8gAXVkbB9+CVRL45bUz1m722BReJVhWz7Mg6hlc1w3YtH5H87KCA4C1Zi
cnd+1w+/VOXQVBUHYsJYp/CWGyE/4jW5qkunpzFF29Dxgz35YZQHEF3+JIgMKJNmX4tU6+M4efGV
Ye5SqGyR5dUTvRrgOfwGBOhY107Eo9MHq22msvJt+mTJqEiVQ4ls7gwicNzK4VkVFygg5DBI0N2C
wAoci1NBMRduOXWNpSyYUjKQ3KnJ7bnFnWOD7+ZMeOHJNJ8rYgoM3nbfOA1eOKNjQaN0FnLKfsLf
mYSt6brmeVFWl5Kb7bJgDtRqQ5+O1r6nbMRrm1f8JbiVBmPm1BuyCCBSkjH2gzxqXpCy3+TWtkAf
euPjK3KyDZTdxXjrb5Xn0GE5y2IosLWrqFWrHxWryUw05CCcIqWUrQ9USnt+u1ZQ4131DdvmwEJm
urLM4gbxxxTTtymvQMpWX2zT8ohEb3oyg0hZSe/eoVt5Vbg1rju72u5wKBnpqza1xJAbaxsRPAp/
Yqn2NV7AIAtxChMs6Z/854c3kvYh06UI9/ZY7MlWiOgSZyPIXXCxaiC5VnkyYxJhAFBmtt5cf2Z7
oMtoJNBj98R2KhTAf6U+kV86BSEQtk17VvjwK6M3KAjAXRbDwgMexEz6feR2W1+ZRpc08sirBYoV
KKbRiZw9I9NURi3CUaZ5CLLoNmUBFdVOUPTRMTsLeZuqjNznePO2KQRY2cqJTfcSBT02W9jXYyVE
IZu0Mz9uVajHa/scjyjHUQsI8bxrMjYn5ZiRliSSzeoXJP+ga3aJZ8A5uWpvb4kc/24We2r0uOI3
7+wT1Pt7yS6QQ/zhxvFchwbbwp3pDOjb6KNKRE5+q3SZcACnDgxw2mF2GlkmyvvGVMPwhT9cRbRL
4gkoyQIMWV8F/U2xs+M0fLkV5Eg9v7oWDvVcWUkhzhkzKw4vrqKv7ZSzPNgfmCaf6m3sJv1y1BWC
kQrB1znrQ+tp2jWnLeOZjyHyJVH0on0hdpWJrIdLdpZZHmj580UZ0I4hO92lxPs1xPSoMFPx7YDh
0Da9Lp/YSIq6C24uhFCU+mUirXGFErrhcz7rrjJPQOcTSe2lAdgECfb7cFaZH1jrvtMfx+JnOU1S
E4hJZXU5VVvuCPeq746UceDUiawOhq14HuIlM7THSIGxJyagJbkJn+eXV7TFdnaueK2Ao3UYQaRa
B5NMqyzx1aCiCHlpIggQ0Dd4HirzLDHO/R1ujpJh5gaAT1e8VVEIvqgLk0NnISpAgjZPO5SDW6Qc
O203RZqDF1+LQp0hJrFVP7FsMjgCTKw0sCVHHkvNPo4yswyMcgE5XK+4m8ELU4LJvzYS0O6FQV9j
nvmciCrnr8Z76QkJvIwq09krmNLlNqaMcngsnkM2W3LIOafOJA97oTqudwmLRkdtTG2d9uUSITjK
D1YeObmLUsqDXt90MSC9Pl+MlqDeoOHKxCZRhnJDA1d9xI54YhhU7IGkZToF5uuV7NVgO1GZng6U
Ostui+3MokRskn3b10mf+ni6jqyZMB+snd6jkbNa/hPIodH6LUJXZjyEWv9V9av/5MdwP00lh81o
0Kfsll2lgTmXeVjYp7O2JDSRAJ+zkFEbwQaKYbEcczIpo8/I/VNv60A0Nz0NY3CBlxs1RSsTh1KI
q2DT8dGnRCOCC9y7tipuLUBNQyHh79NCztMGE9p0NBS7WExLbzKABzGBZrxJwQ7W/PO4W+uwhpTb
heJ/r5ts+6hPwAo/JwShHK2YBI7EHKQk50SYpCZx5U4TIO4xLeqyoM9fPXGUViGXDqpJ/8yEQiHa
tm4PcQShqWdPB0Z0tJqFHwt3+SrwdS6WwaxgAc1vSj+nuVfIcGUY3th89GIXTiceos/BBYj0ff6P
5bWvYl5aMrVCS777D7MNWs4UzUSlSfI9I3a4dD9z8mpg7t05mh89e+OpPI2PLMONAyW8WpBCOeCq
vXgAn5C7zukwD1L9jWtLDTUTl07IXJCrYla6VgXuhR7YlVVAyQwUhWdh27CMugD6FcELn+DdbxlI
tNWHijgiY4dJ0ss1Cf59ZleSN2hAsXYOcAHWrdquIG0hJWuNZqLIU5HGkC7YpFx20QOSS5xDiCzv
ZiHFPxXcbTx7K9h00/LsrLwX8Tj/XeXu8oGaMuw9ke2jZx/VbxYc95Tjo9DOL8znOoWzXj6azeGD
0DhH0CJwCnwbFcjcBOlfsGl1n+sGKDYutrNJTOfh1n9NQN2U5/cFYfb7UAxUXhaYtVzTq2FPuFEm
wbroOwFhPLS24vvm6NzEjztfiFxNPRtMIgB8FrV42ktUvWqdaPppu3W6SMi1O1KPfjZOwpncvyJD
tFVb5G+9erBfSpXbikmRVbvCpgVo7dnS/v/Y7vOPZlaBgIOLW3yu5FALCPyT6v4UnLA/5MPoIDBu
NqkN5hB02IWAkPORQzkyrPJb9XE10tVrjMmTMphQtMn3QhzttSCwR/S9Ntpbiz9nIcMefTlGF6pY
2mywnFyE89T/qbO+hrkUb7YignSocSv8/4bYlNEzKd3ekBgjnrfyrZLd2Z+Xc06kJ1ppOMkUof3T
ceNOs6pcCWcZLvhp0cbM2b3A6TkVhbWeivqdV1Y5XmHoKK97OsijolLLbT6Q5e1K3SbUlB7S0opf
qToHZD0bV7LlkPXBf49UbU5rZ4CuQ3aX24x5T4F6X6ieFu8Nz02HYYXp7JbnRx8LwDMUTaoo++fx
997SH040jB4ozPluzoKhCr4/5CzaFJM/OXRx5U+0E8BZwZE3l5f+v00QZRZ+7sv0pg1BwK6zEMrx
CwdnQN4rrwEboq62NhOTOLcZcaGnT/wtNIV80jn7AvJopzB7kWRuexVf4mMa12vJjtcqJBNsAKTk
QyX8/I2E9DZjhyNsyEEQubSiUWe79d/kh3kan2+HZhXJwK5KTU/jeDmqPvRkJGOk3rmmH3ZQLXzT
5sR8b5QCfFvX2veCBvSNfdH8wqUWa46Pph5+rxv6Sa9Na3xj/XY1DB6N4p/jYOUjoTqhiE5vq5Y1
jDa9NHjGhlexVwvRyAH4H539XaXfKiH2fzS4iCxaIrFE/ecSHXzhIgBbSvY2UpaM500BxJSrSGJU
tltdYTzy88uuyu5Lx1flu9UnYEYcUXYbuzj8JI1j4scYy8qUNSKa59jNk0qrsbVfosd93YoxINE2
Me05X7xYciT8Knwv9WDh0M8JBBYkwSJk7CrWBfk733I43+9Hy6LIEOjmF6AiHeeEn44lYii6UJQ0
TV1ezqtl0UKgHe8SbGk/lBoCFoCMN6JrxgkC6P7oMGWC4O+/KBhwRSkD3k5Mk9mIGC2bp4+UY5mM
fpq0DWIq9Le9YI1Ru8hmV7a26dgXc7WLGysUwSgaFhM8DuITSyxukoXt4W2hy524MD9zvPTQMhh2
O6QuYBCbSoZ27rLl33DJEYsdUn9E2GgSVaV30UUzHjsNfo72Vy+jRPhXTtXQf5iNZtwyuR7175zi
NvOSdQS7hwXS+KDunEUvknXB8NE5Q/0mBWKKYQr/h4EOHSJgreQSfupSEhzvT/yWiRR8Z15XXwar
Mp1UJMI0CK8HA+pPrSms63ylYqBUESCvZX88bhopD/pieIQh6Gsde28Y4/yWVx5O/MUOXejoY4SN
S43qfaDg5ZU9HfP13OFlRhzs/V48jGHmQX6CpLYF/Q10RQxlrsR3oWvXCp10Rpzh5ukyO/EenBji
wTxy/zg/Yg9fsDpZY9MMP4fAd/SJOBWFtCPMWgPWhxQmQFJaxtm/+NpMccVNCLgwWfH7XVsk/uek
MhAHTtD/apVM1+hBn/2cQoxWacezVE8HDgUbv+gX9S1dR4YqeKFceP6klry8/wcQ9a4Qd1hr5it0
Gkv3q+inPRhFWZNzbU+Hi/VEHc2YEpsz5hv16fGRQkj3SzwKKU657JO8qxXwVglyRw2BHyAl1Rn5
kvplp4T04YMWqQi47c8SHyzBxHOJ3WeoqLrKxD2SyyoTR5lyBiEIH/Ct4bmjw2xz0DTRrSDkGzVO
FZL3kdxa8df/rFO/i02FqQ+kRc70P16Rbc+Fr0HKgzR1NczJkK2MLiv55pgLG4GfMSzveDIvW3SM
IApAB2SR3+xObUdYazLm3/VhL/zG4t75P43Qt+F3fbzJkQ5AcfBXi+k7dvpym0GMbZ2L16gAIcjy
MTdh3ExRRp+kK7H449/j6qqL0jxO7BZO0stHvj5DZZf1qY8akRJ+HRBOh9tdGsJMLODLUZShTJhu
iWNhjRRzzbDBxwzvlV5oZMHm+iwfjLJK6FWW8kpEePm22hBChHRfO/EBMXbdwJ+9PAz/afargE6S
7kHLLQB1EMX/PdzFShDCG2XXctkHMny1uVkD5SI70qB1sDQ3Ks8DDXf4BSEX/2wuAwEb8oH5DxR2
NXwtY5Jz0lbm0AX0lWwRfVGQxQwa4bG22Me15MpzfmskHLfPgRI0cjnRIlPNq1ZFldpF6UziNVoP
/95NxVUuN7LQ2aKdJ5KLg39eQ9TC5zMfkTJJekJ0WatVPdUhb3b7Y3lBENrZHQ8QkKUVBR8mVVnM
9KiARxDxmIyFoDpiwFq0fswaaqcO0a3nB935cJFx/lveGBIOj78jwTa8/9JFgXBi3TbellfNnyFz
ZRb40ryOEmiT9hIXN+III5KdjSYFHNekz/6YyjuwC6PS45kswQ2G2Fv8kFf+CWzCpwxOGWVcSUnF
wRYl12AFktXIwE/lFrAASLb55XcjiyKvh6Nqrud/UPYXDpdlwLveLQqjWs7TKj6Lsp9PoT4F0jRb
AE8+FzlmO0tJPZVY1Jf2nTy0guARPWH8wMBc/2qmwtua13W8NvtP50mHowtPi+/OlX2JhrJPAWVo
cxJFj7h+7E+qweo+F0AeSIBe/Av1rCaMxFupsUdX4Sie6tz/fKk/VuvnVQfhbwJOnEl2iEWXECQM
a7R0PykAGvN2EPvEWq6ZgUi1Y0sh9T956frv5oP4w28qdc76HBYNiRYwdX+GK6yS4wEiz2Vdvh8u
PjxQAiTz04fitQLqEe3PtWfiaEDbGzSC6NL9EAYdW2guIp4TBHjjwVkfvy/bBmpE01Ttfb18kZzU
VpLivDkBLhR1hjjo1n+c9y2DC2g9SS6PPL6TvDqVDm0mfXYdaEBkQGp14c98BuUM8M9dZUWP4q13
bw0q5ISgvJg4CVFVYo+EnQSlFpPTII2IrdwNQZqk3grje5PH9CXralN3F2KTdXRF9x1oKAnReYr3
qYMUew3ElHmunQfY18+z/Sn9GSDLrI5TlxGUOmGDwwA3UUo1CmdO1Esut5eJvCr4qztAzAsZtOp2
Yp/frfUToqcQfYAdojLqMPHGPlUrHoJvBYk2Z/ZrTXyz3jqF4u+gByiJ6Ccg0zrJRFjmVpYbxbEA
rjb/nYirlAyn79WByQyQ0hqnpFEhVS/cj6RdfIXgQZMhmFZ2Tzp7kCJEkFmBKGG4lqLQeZFTKKFe
pK1E0va5d7ceUZxAA2VNUwlta0Edo+MX8VPhWHCeq+2/Drf3M7C3ZHDes0kd5y46o0YeHK2a1Ttm
jrkLmpflX6h+ZaocnRyfFN8v6RfcF9YWLZ3ChLhjHVhTYliK68Ag8AZi2/+ISjaIRova+DdHQ2Pu
Kxaq2oRzZQorFDc3lBQz340dTNToUFktNrvBUNP/Lds7hWKwjrr26I6o1ZH36xaLn4/uKymAi6LJ
1zVuZkFVXr+3xXZKfLwOqq+IMv0ju84O6iBWdxOxqfVj45f2CP0baRqX8fORWqo4m7LiNR4kZLQY
DGW/0G5wulvHonjq5yoocdyKBciyeR0fqMmN6lGiYZirtUqFahCaZhaG47qSYg6naRm+BDpREH22
rHHS+4SI0OcWzalF0QNN4o1Hz0tUYHWJIwEf5rS1n71DOtBzm6K1WIVOJU/MsgelZedb7PhNaWu7
lBLXpgZCJSpoh4HyKxS+5kzoByIu5X7ucBcfMJksxkcYzd2KRQe+oVuLS6OayicwhR17I/g/DzLq
pmLPUujsycgw77hF9a4dwwSjFCUyEJDST6F823YU4AWyu/mFBIrHs0h+HCgZoveFBQhKj917Eo5f
9tinrdqcRIxWgOgmp1JwESwhjzZyf9TP2aLBqvtDgg4JCkvbUICYPDjKqr/fMfaHfMOwdLuAdkuh
qXpbGZHggRntmcknW8jMfS2hGCSg/VGemhG1Ci8pqQB+PoQvR2012dD7hQjtl45poKTcVbZuUZm8
xhzZzL5sk14xNY/FsuQUyOdx5bAemEojJzvW3NnTcnEDt3wT3+apCjPc5Cifhj74WQBUIVv2jPJE
P9Tt7mTr8h+sMWOZWEEhSPun6Qk1KSiqGbD8W+E0rprJbpYUawxWMZ+sHdurHQQd+0znnNa9ZpnS
Lb3iWoFplS6NaEuzlF6+dtUoTK0XPxHpcg0cHlauRue2ygOKbV6Fp9Del8Iel6i1JN0838Vlz/P4
B9SRVI2x/U+Qgh5BejKk8g/VBRKkTtUsuyalvouYCPNjTNZ8QTBULP8wxUWZOkb4uoHHPlwgc4z0
Ja3rkePnTmpXqMY7XoBysY2tgaGdQo5/9xi/0qmuqEHeCBtKRyQaL1ApILpMbGqxEcxprzM1m7hZ
WGP+ofDTANmYBj5ZUUTWFYZOd+rZZ5bYPZVMMYFlaTXb4FiO5boX0hWKswnJgR7OUrWj+s1e5bdy
vkn0QrvgnBDA7rYdhoEBqUnTwBfmeKs5dyU68TqnOzkSLB5V5B/66fsn7/19iCAU7CfbaJKxfpq3
OVOcJmfpaj5TGaCW4OCykKEbX6ZJi/Fm9iT5L/XpdWFV3eyFaaRBTgzwZm3vwdQd7XiOBcG8qMkh
9D3tfZFX6yeJsUlx0BY1l3OuiNZ0EXIh61sEZsd3yJWiii4cEniosEz2bw/aljci/MJT31Wy+8bm
3urL7gPTu2Q5HrL7ZIWnDD75Pkg2EmoY2QEwtUNDRm9QI15jO3tuXN/xt2+f/8bTtuuXNRV8FdvD
4yzCmxz+72O1UqnGsrRJVl0oJQM9tmcs3FyV6FtFvWI7f2ZZRfqOB9Lh49XPUJRv8zU6CPxa07sa
wO4II8V2G08upDmwX391nisVq0KfIRuvYNPoauyUkv7JXTuzpEf5qH2pA/qWhFGpSVMWs68skMvO
dSJAfHbBCwdBIksPM1PUACRrmFBgAyGm6IDFK/vKDYIR1izFVSLdRtoI2WJLKAOWdlnOU5Fki5G1
Rommd7f3nGJDqNx4VsDHIcs7aFtaD325cV/ITzQSoHeNqc2ygEBhbGv6ps+lRZBjFPbuwFuMZXgn
oNCCq5o9LKK9cCc+qJiNHGL8S9Neu93aGYvUcvhqYlJTSdnenCn6j7vXRtunf0mMWTMAId9dMYjZ
UA7AfOK8GvDGoTde6LG/0779CDsWGXcnnKRIRyzUoS/TZara1D8ib239uV9ScdbFMbtrgHrYvlfw
wysT4uanEcU9q9TpkW/9hH+YX0h7nFi9G26qQ7EQoXbRHViBEyGn1cInYjNIAGu/U03GUNdoaO9c
v3TjNhmUOQxuFjVFZj3Td/BD9QiAzKwJNMZvShXDhVisOqa0qZz2q05iyW3RPELB94/wJYRLw3G6
7xUbf+wCcPHrcr+FJ++6x5lP9dHNf2bC+/Td5umbw54LrXh72TWKXFNHzXphGSgrL0dz0Brz1+AR
4CZCt2E/LJHmUxsP9tf8U07HReNru/b1lu8eRLpKC5qaSltZJgZ9R+WfZc6G1EzB1ogjJbIaL6TJ
Ek8ycEkAN8itpvgdpdF1wKsZAGC1KKQRJQLWPQHSNFCJnBokONSlEpFJkzMLXthjy8+ZTVpKmXok
FYs63JDqZxql2C49xtTMOAqo/njg8GC7Y6OtuKwu/U3/2z7ct+/on0ByLDVLXvimW9Isp8pD4xC8
NAnIt7Ha/A+3lqhJvNtwQrtAezftB+mlCFJcE0+w20LTzQM4HgbhY6v+0qzZjYGyPllDlvZzVUN1
KkrnWESb+4xHpEQvzEIJ0YA9QdlOLQauDQFbvQrj/aiwiFxGdF5gDQNj2IHCUJLXcxeyIkq2Cg4G
xooy8/GP4agfM0V8jQWBbr2ZvuArsNIL2W3qC8YL4H+n1wUWg+ugMTgotl2NVZTJnN67W9hjo04J
4gwvIyLp0SXkDLIqof7Z0MivaIe6BkQxRmvSqngj7gYMGTHDjqwEGNXC1rqzIa6osgVKgHqIMjzA
Ynm2IGw8FJY++Vb0QNJWGb0sljtt0Y6vNT9FSYaktiTOa25VnQOehNLncqHRO1LozKrivamJRnQZ
2l42xAUbGUj0xZvch5RA+AYqESNN51xtetpOWP0gPINjF+u9OMXZ5MLy1VZoe5+JCddWz+J7DCSr
zO69tdoPJrJNtZSC9aVzbWim90lsZKETcbTqE/Hczwn8iQs60UtvCYIZDS5jS1YxYrnq6UY95Edw
1Wx9eD06fM1Sq+nRepazJC1JQ9GOFdB64kmjabqLomHv2zQK5GG3uNWm9TQmkNddDWz4DTD9QdjX
QbSYqAkUpRtH5o+pUdYYxqecO0wzZIwMn4/OBI6n3R6K3oQ01NR3GWRWRthq+okg432yPuE1r7c2
C6B3Ajlpq425Wncv7XutVwqr1oWei71yNhHX/68FzdghaYJ0s4cHqNiHb28ibTvqu8WRXpuKaz7n
24GeokAj5w5hqC0iweedgkclV4qwJ2JAulliOw+a1tJcD/EUYBxrofPpGnQopiBDAE2Q0tVHzt4q
DqfmrsLfUwPfED8/AJDCPln36VwcKLTCPoFDcjbqKCof9VfKx9AKUwUJ7xDZH0EcastBgNYmcVHo
Bg/+bYJUeynh281Tso0iAx+gd0KHK0ozmTHynqAXrFYuXBOg6Wj4Inc0KaPGg3NX/si80ggk2h3M
vGnqidmlHARMpEKfKKHqdd/LX8r1pKOvWNVVVEr7e2KlWs5Y2rGlvrDc8NVyZ4EqllS7RvMvWE7n
eFeY8yd81AtEmu+yjIlgtVrXabRCF89Cvliypu6xhH33BYqJMp4tLl7nCSJ4/X9EBTyKcPFhcEoV
3Z2mEsy4vCRfl8MhDZ12KITJMx4txAg8TBp67VG1hLWaXF0QSOsTt9OePugZ5C2QPVaKCsobnekU
Vi91ak7mAawoLKXHyQX5gakItDIbUkOlZ2H8hU/p6pkowDzYugu+AQLo2ChFAeR1KeZ1BRV4VzGG
i2lMhlO9vVF/6MMRLr+H2Pp18rMRL4Z6qt5M3FHztiPNLOtMxHzQdAvXvUPDZfh+OD8X+kY5/1l9
Fy31cg2P+5FOhXSnnWVOXRUSeDH4H4stoB/1souHPEVTDFtKEbqnLdFPDC5vxnXSiA97yK1KdRw4
8AaFVVtLMcGuD4wu3EQkS3sek2azQq+0hjKxwVU6TjaZfLDsI6+/oYL2HdVXgqkizjTIwjlTSYTV
qRmlCunNdT7/mQWNviL2ZTzEO6MxOH7BTX+becVAEHmJZexNC7wszjzIfhUU4evz1zykF8EIvIT5
AIOSqgWOoH4m2QBPsbJ5+r5YBj617YYS+jAxNXeL/RnZQhAqeGOpwuENMTWX7gtecep8/LVOVPtZ
3FhMxVVo9AOjxf13l8olzuAteB/r5J+ynGtr9rKzSI2vkXu4sxPXQiXnYexuP1HNSreOiDXjU6Lb
ma9k/tKKgs6HqbY3oc7hMmO17HRIs7b5LF0Wq99mSkT1h5fgPGkFqSv/MmRC+Gzm8tuUxpnTkHZM
zLZzyJjzdEboCL+3g3XAMWqmOiLeamfj79kLKemGtaseJdoZ9Wkq5mGczpcRDD/y8VaBNfdKKFkX
WI+t8KD3l1Bs4i2CJUPcy+mOmCGQHf5R7WdwKE3DnTt5wQsGqZhn2Bu4Qmt/Yiv5UdHLd6ZQ5BBf
C9Cagwc2WmGfAXx6EQ79ERxMXSEqls8LDGCZ3f9t5LjT4R6TSE82nri8zPf3hMrtLpSZLwhhxs8J
qpd+4dK2F5upw9S+nccz/92j6hL8gbE+962vZsvVVIxdPKstx/Ns9/AV5NpVsz0tbiuhW11/6KaM
NNVRORZN9FJD2StCKDLGvnCIjW5FvgrJZMY0H7U8U7Sp0KvNdRYSNw8lwZJGL/z4RHZe/hemxIdX
BIl4fNk7EySIuIERqB7iZD/8Qg7CBnY6BdObe6En5RgriNxhQNcuXrdi1T2t03uI0CR8z6aXc5c5
LQL30lTrLAI5G75QbvDLqAQexF84XezAKljMVFuif8zXpylGvKYrEa9kFS2GqZ3cJ5GCOWrCZPRf
xkbo1nOEELAlfgLdRH1VhceJ6nwq6ZXni96NrKhbD/GOLqY0ESTetjv/iV1GMp5va7XBfQguo8fx
vSQ8zy01vw0t/jwmkif/jrPvwyebUq+4y27MBR8yzIAnOf39QApOPvJr+0OkHPc8Hm6TtkMBH6Gh
BzULHfzoor4eikLaAMfUAFVejwsNkIGws9XF0bub7dL9nfR8IJ8lKR15W2XenNMLssMkR2A+K5zh
MGq4qA8Lj27aQ4P9NqKhbQN7e4+DEkD6DGLBJLOryHozxsVBi9nOueME8vzn8G9Ne9JjlW9SJDx7
gjMEMYwAJltTDvfnFaO2Xdir01L5cV8DnqEkb18D5cI1ccTkW2uPLR5VUTY4Y59M+HoAvzZbN7Kc
Ww126m61oEcl/RNTh9YiMmksdf6H/XlmVFYXzZPPWQ/Gz3Q0HEl4UfISCDklutpFRmw8cuMQ9GMt
UndpaEElke7IjLDP10YdqtwTHHMP0yrs62we+mIjbhA0fvZoolKXJiOHeyKHb4AdyWzUmBCxc5Qt
i24ILdrZyRxaHJh5WqsNWshASge3ukU2ZhVmBNyisStWG7fRaoKnnKCBGULu6tcqmVKbese0tNi0
l/jRyKs8JCVf1U6GMd67oKZbOO/ieoDR98Wm8UzOZunnjDlAzPTK2qcxHUntBb2IbrNT0jowcDKj
k/bcb4TPAhl4WKxN/VnJN0jBA25yZHPJE+Dpksn5vAKFzEQVebWBqLAeH/GqSKVdJoHCSHF6hVwZ
+NXBdMl+lTnHaHG1rR2hkb+tjnfcxonjHOiuP9GQJnbyTdyTAWGmDv3MFeYpZLzP3QpLN1Y8KQHl
5NHPVoIOjRVQ/5RWIYMjZ5GHvAyg4K3UwarqGR/lxSukzUVYsG5J/QEfCugBd0bz+QQ2Jlx5JQp5
Y3VOUIQmmW7FfrxRj+gMRI30CTAB9aAN7ccYWOp1I3urR3qy1TGNxCFBFdrxq9wx1s60X8jVryDG
oectzff1kSN44vVJwmEzxd4AZmqXtoAlY1HBInJ7kgog3HUOjLVE31hPiBW1hG2cDfkCwWoRRdoJ
X1O5J1wn+1ExYzreRqfzWee6BVxUh8WVP5PGhbZ0QTmGND/DZsGmMT6KGi127AMOEdXKLbZLE1hs
Jl1sLQPeU8pLe8FU73GSSEjfwi/pERx62LWxNRQdw1q7L81Q53UGjhAYUv9vCNc9KLyn4EI4gHM8
2qhRwjS2H5LQoNAtF8E0/d1zKdMiBIoXkySYMIkXKYa5QUSeqlJ4bIq2ngqeL+PtSnUbO51SIPhk
Vm6NDAwacT6g0RGFtvpaN5RWNg0vEvc1wHsurWUgT93lyrG7HiBbZlBbRXnrah5FBACBCzAmPUvf
DJF/u3wMVpnJ3gAIf6H7pF4N1Q68cJdi22gHN78N9aYip1RE/gOLrd25yLe7mI871xSd3tcdsN7g
7CB78mw/mug6v/psz7XkwhnMtOZ/jOTSLU3SGN4SDSkJAatSaTB8WY2VmiV4253hDqbZJhQ0RKTb
VzwB79aWOe6b5RCD/azqvcMczbizPePuobQf8fpE+/IpM8891wyipkEI/YhKzSSUkFvuAyuEO7LI
v++BIyZsLu3q6fOIWrVgBOSmkaMZJ5Z3GyqXR6z86CNTUqmVd3AN8I8TvhM1TwTp7kx5A5RVLcNG
Is8xMprybkHxxE9fT/pZFu4fuokBywxDSOOphjRYlabNSx10r9SU7NSH8cinkUdUF/d61W4FgOZJ
eSFPAaot+q5lldtQqLKrYIL9TRfO/X2tSsfw9em/iex6ijc1f2m9g6FEpPDBMfM8y37ytipN6N1Z
XJhWw5OT5DIp9se1x9Xe1EOcU3fibSFww5be5lnYB3aj1R4LyBY7Rh6kAQ/wBMqEOhwJmjE+Fxlh
OKb/hklK3ufnSe2dREJsfrTI/OMze/dJNQBxz7/8XPwFuJo1cpLWKkooTqmio7vJLR9pytaaPeZa
RaLoQQKlItc+kq2+Q8Qaby314MT4u7GrfkC7UU/mq9dW7DYIF+70I5LKoyln0zWe9RvcviYMVML+
+XYJf5wlK9s68ouyThX0NhONXb6mXeDARie1xQVr6i0aiX0E8JrAZGmZzBx1xYAyX0dxch9SCX4j
/nAa7D9Z6vcfX7yCsf+AKriMyaLsgiZ+hi7e+4xVdvUQ5J5cxbtd56J8Yg/bn/PSj8mmPBUvAVkE
apC09P1SV9YF009EYo111q8hPxh3Jhuez+28EPmUkg+25DuSzpy80xflV0HR3Fkw5WSnxSi7lKI2
KQce9qPOZO3GSzibluvm2WHMRub9DRrMULGnt8bk+pMFRHdfY4xG8zO7PiNzx1x3zFfCUeMRTSe0
+L7IEmyvWZITlzKrjHV8JibfYexJZ08cWjCTrrFIAPLw3qjJE/C6NMYRtm5KWTe6kaQfXmMjSvin
WNlIb6opeMP+nUpm0lv3x17BMV0owoMyBqvcZwR9FTiEREEZYHFyXDpFcImsJEOyfB9+D2i6TYLO
wrMPReyw2ijob4LwM8GOXz1Bub1aNbesmlmtvPLUlFlwvriWgDf6pLgeb5AjrwRUdZZPLg+WsuJX
iTOys+x1QEe/jui+SF7NH/PQaBmca1q4zeQUE0AuXsNJz1HPvAgnW+eFS5+Lp/BiwNP9eOpuJmqF
j0UdoyF0i4UVz3aDZaxDC5xXhq1KrrYXiUEdFo+ahalTiYYbY0ejC/0DXSWVLAsVwwnnDPwd9V/k
SKcx26o7RgzEpp7OgDDL21Ghn2IxIamML2F/D2zFnqzE+fmtdfX1lAhzOD9jaeCNLM6XCVry1aKl
ZETsriyQsiWnkTM+sWSxhk7KxGu0fInB4JUJCiIYg3Y9FWZF68TnE/MviTtalV6VsJW9PqRMWZuT
ZeLO1ZSMkr09wadBrtTQJImGbZvY2f54ETh18nw9NhbbBfNiSoQlZ5RTAmCkf7kYIjAs45UWNITb
K1/LHKxrdiylVMBAqnU4LOT8gvVhB0HJPsP+mkGqv3EUUeKVaT/DTM/y8L8Z97GT32hRJn1CurFf
hQ6b1NrXH76TWyNaWihySylFO1BXuUDtbevZDoynNetJADXCQd1J29KeGe01kSsBXkofhGA7a8J+
oxI5TSuDJnJfAZpK8TZsGCjPJjiidz/oG+6bBCk/IJODxw6iRsBYKDcjey3xMleb/2IkcF7jXlLC
4OVBi1k8tHgBB5DZ50z0qnr996Ml0/e2gsljdhRMspXbUOW+sc+QdgrHCLzk60N2YejMdWYecxEF
SBBLJGH6183YgbHODWHYBogl3mo/kdjd7LNfnbUOyDslcTpQoUPfjVbOQVTzdoQKcnOkHm7sd4aM
CMZQopXokTmY0CLe88MsztmvUqATannp8NrXcgW3ZL5wtcHs+umB4WJLbh9ZR6nLBdT8v1w3tSGJ
NHVGBqezF+VmXJBXEqUcOBiPv5FtLliH4JcPqw1cSQuZbF9fGTfHi1AytGRwd9PJ0iNNJt3Hs2E3
3eraGddibaHbYk1Ob/m29jcnp5ONgbxv6YiedMV/1aYYXDD6jLoZThfKrCHxLJN5VJjSwhdIhY23
V4nzm0yr8T6En1XTOTOJPCWmxhc4NK7580Qix0I5qkxEOKcSLPPMk3sT11rM2XAXozMcvfUxxrva
ViUpTNjRDEdld6Q1NIlohDKeoKMFdvohDjIhVfQQ7exkqjYMg1SmH2iOfI9CnVp3q5C2cz+4MyNb
i6dKFqkvxCK8vu2BRigfi8ylGD2+46Vp1MMpONNNiU4k8sLVk6/c0IODywPVms+Zktg9LRGVHdta
RmzedCVHwiIuyYuSt0YxeQKPPuqtkfO05mKQB7fE47BXtbcJWiKYYVBz+byZWvMmCvaXrL2WWz3/
OhkITvp+Ukw91Zmisqjv+xqnN7uBO4ebDAjUC6aVpkyS3CMnTNJ4Aod5FmqZ6O7sfWo3lX2Yw2gO
N6GU7P/hLNLmF7RGwCajCfktJI/iqMzwKy3iCdRiSUYdCJ+bl4+L4HyTHH7J8TrvPoyfdtdkJMO4
qZwyueslNiQ4v6nw0iRCW6kcY7R8LePfhOh1Rj25DIlIyUWDED5xepc2EzmWbyUN7yAUKKqyEjMV
SI6fkXQ/uZqy2Hnej86PAgRjLit2CxjlkPHkP6s/sJqenaSelMpAZWrW5TjJxGC2ODg1cDafb50q
3IX/c82GGWPKSB/mBaDyCYf1eNQ5EHm5cvt3u1JBbD8CeXoUP0zXe9XWDY3Zn+6rAiH5lVENwN3v
zYcodVfmQ77+D0rISgqPOYMyvFNcqPYQN7qCsejH3QrZjjt4bwW6LHQMOtqpG+fZYp8VB00DaSso
tE7I9HGOzGKTROG5/nIaPnTq61p38pLpnzBSX+6GVK0Htfmf3YGUEyXD2U3iSY5s5aQWWzWEkIj3
+e+sWjI/bHrtcU1GnCJHbdjUL3qqwYlZx4Jele5/3lqCUyYvdrDYedTK4XiFDdJ0biv+sSeYHury
Ynekuf2wlyCVYM/36zaZt43SCtePRLoOy8oSp7Wf3+mrF/Lf6G0XaL3mS3uZvrGVO6ANGpBrgNEK
ZJQvqYDPdnZZYQ4ElGc+wMOkUYkXJVcu6+fEubCIsZrVRJFmoj/QqYYrA0NkRQJP8HV3nthjnhyF
2AL9TEfCCMHNqHyVpnG8HjgiXq7i/C9FnNgn2VdmwKrM8HV0bsnPyQvYXrEoqDh2BBJ0au2vjI0h
Rl9mZeuku8rI146OEzBT+swHjW+7z5uI7d8aniLsCDijMi4f4u/ySo6aYzkqJTlFY5t05lDsIWdY
KkLhHkSOT/5zKOp5z/+3iLG3oGR43pPGiaf0jWIvgN3Tir6br3T5MziuYMiGNSNzL7EOWp5whilZ
aLpfEDKykbQNSJMTOL3sFPTHGjvD78JibgRg8//6etB3umbgtr2Y0hcyyVqbgYPy14MrHNlb4T5d
Wxir2bXWfgSOYvqelXNj4OJbrXzuOXwHuj/pxddHDS3MCmjYEDsdCn0O3ynYeY5GS8iLlRaCCR7f
Ew5jioxwFn1uZgQNB5TVET+wkxpNxZIyArJF8S7ovbbrDnrCy/Yf27v5ZtdmYekUdbLvRjkwxicO
HWKy0p6nKD1Nzq+jlnmjpl1TB2w66gl6tVwedhp7bltE84UfmwBJjefmkMYOtZGry8FCC3SWdJgb
ryfmpvEBA55w6DOS9NcaBEmwPZGK0L8FQBwT2qrWa+RxcUa6IbQ7flm1jv+X29CrbM4pAH94EBoY
+KmBpDpbXQGxjegG0cEmb0RYvaoUMXbjGuWXwmph4D/gmsOSQRLYlIOIns7GvLEN4cRoXVbLwcQV
ZSYmGilrfs0MBuGpcpPwLZBI6sA8gdRu7/UGnxXrKWOoEPFtoh//MxByoSUp3LRiMX+2YzFdT6a9
V4PKUzEd75aocqXj1tYSfjRfunPTE1WpEfZXdN5WxvUSotgK+pf0sO/ULt9QiHf4ELyoYrk+lfnv
Psbadg8TPcZNup7qk8TsD6JS5XO8EAAu42ako8BD4AsMkvri8ZBwDwjHe9I6xeg54BaPk0nEWaBc
G6usAis4o6V9aAXE5UXgoI8mWgzQpMvlpmzNTme79AUu7GqztJevd0tevuuuhX3LGKN5PboMxkRz
/Dtx1O/lUImyQrY19sOnXM3XzGiBJ2UHnvkFxyLbMiA4NGLJHFV5NnBnoqTSL1n8BIPlcDTeARZ1
MI4nnIg06eNaKAOVKtUcaljPJEVlNvNBFA6AtWqL0QoImiwxVEj1HXZ20H5fRdGXHpeRNAOdc1Gj
s7ExnjlzmrXMRfxrFGd/kOPcvjS6lt5u4tQf+ARmrY+7qfvu/rKfIjwxf+u+n7Ukgx6qSIHuIGGO
iAgUffDiIx+4dPKds7+/G7+nWzOUKFVpPRZ67gbOjSHFaLOaAK5GXLBxGkDIlbqgHjvLK4/OF7+N
vDcOZHYOzCRqEtJ8rr0o8DhHRPFbFHrZ5rdZ8vg/ykk4YFE+SLcwQEJn7YGltjXrPSoGNo7mxZtJ
g5jHjuoHYkJ1dDFn+BvGJahXoAWNTYspcgQGJaWjYyorr8Q8b7GOiEGn/5/sVBCxz2ifowcjj7BQ
Slfk9Y6JY8XryYUwLFKzPmhl2Tcy9CUOROlrIeUuK7pbRIqfNwTyeS6JWdjyTgIuRqdkjeEtyKV2
K+aUpJJIHwz322fv7mhuDeSbjjHJfOc38WvY8H3wUcri0abVZ+dO5l5FZrHSkxzH3JGVl4zNjFgK
OzeBpxcrKsHWZ/nwBxj6vi0QkHQYEqtwZxDTktvUTqEdTCQ9Zx+gMl1eI1KCgwAcJu17RSVzpb3G
3VUPBEdY2YktEHIClIu5oe0Mro/Y7KhzNHW9QLTS8fTo/w0z94zBlSRRvEP+DwQOh1Xb+rxIDlDB
hUNVQf7b6Bkitv+wJ43te1bR7U2WCV+yCxUUKRSWKqNzO5oZXtPHy4ddnZeQRxVelqbaBx82oYeL
4UI7iNL/SFnSIkRVGjeuH3W8Z6G5RNgKml1VGzM/gZrSdrf5MzyrX9tfurMqHbF+8ii57f7j8QkM
75fwjO2nY7DYEdiWMRgj1oN730LEbkGvZs9cpv9Eo9zXs93ANsaiAJGRyYrq5DhEIjBT9XsY8it/
BjpXNKhjr0Gzew6UexqdsfhayOhfkWnZ52k9opJP7Y39LEgXhqSyDCyc6c+GuYcuQzdWcYbHo3qD
IRtcCTDBeW6VSpVnLNsePwOGM7bvcKfOwrlyTS26Qix/FiGnPTTzAdBJf/vM7croXdLKgqLo4kvq
on6juHpH138Onq397MkXciy/6H9mXbh1llOd3gW/yDCdF/3qMoncfhG2Zw3fmbV5QlfJ1xhoFPXu
qg9OocMRUDo6YhHskwbPdEBd4C9Ekl/te/qbcWsty8+fdrd66eP1A/A1hgPtGpYIZPhavToJBzzC
1uj87iHKRnCT1fulOoB82BjC5iWYQ26/m1+iVlAHdRSNzFOcuwDz+Y/Hq/jeerkD9ssbWxf3ioyV
+tAuWTM4ToEanf1JesjJRXCCL/j+vC7KZcGZAiGckI5m0JWHq4ccGEq+S967wdTFcqyy7zd7mdHZ
6Mj5df12M2JG4mYhX1vlSUbi1yWxeXe974zOWkVjcJa72s9oslJnrbmwZMIpSyxz/AHkm4zoa9Ec
tCfYE9fucUfmC4ioi1cVFtEAVzaJZ8QpiNRk+HGOFRKqGRdG4J0H4zBFKb5yB/Vh1alyekLFtC2k
dSDyn3Ez9ywi2k2Xy7JaYpdJGcvszo5NJR5vDi/8SAyKrdYkRkybn2yrVihXJ6VAnl/FeRTRIVMs
BywEedoSQHqqOcLfnL5L7wloQ7hNqGlnftx2WltLXQ61din/Ahy2EvRpAXOEzNWCntD1MPGeJggJ
VLF1T+l0pHkgZESARy9+TKfhmzMWXvxqfPctQjzh37yzqXSKDpE0apbc0bOQKwSPQnGftw+KHorx
RF76lbkN1GYU1Mg9BtmnXI32vTMQ3lvvqZlv3FGkFI9yYazmyTxvwUG4itFrQB6zOqYbYPgmEgd/
dW1IZrssYsfhowi2jjG1tXdEb2U7NW2b2YntzpUfU7vRxBnPqkxwZT23NF9JsQDf3wrZ4dYEtfgU
ZrF/74brrmfOAnhDGtxvygZqNjfZzavHRGYODDySkZsAUXZnHJqZbdTbhauA8TCEED0vOCOHME2e
eYFCy8Onaqouc0mmHGjyAyBVjd+mvRAc4nhLuvJRoNnHg8lXA1AqNDnfkhzuJp48qMV6qXszY99d
Z1J3bNoKEk7mbuwnFaZYaAEoQZYeL9E9qrYu642r6cERe0Kck9LkCqm2xlbhR5zRfJbJtNFUEwl4
f9zpxiRCEDouqSQZNl4TmF3VYGvWY3V8o5hrH3s6CX6w5U6UBMAR91sDiRhukxYm++w44NpVRid9
76oWUnxKzIUQ3kwLl/UG84szSeZpvcB+KIrGs2GT+eRL5w7/WCAF0FHMtLO5ce77qM2Tsd9w1PZz
7y58G2KbFU463hl+2rFju5Hjmrt5r8prXg4QOJuEB7NQtVl5SEM4bhSpzuYfVKzgfXHOTInenC80
7olP01IRiUJA4zePI4ZMTiJ1ciaSp6o0OorEHWN7iLVaq5RpS5/jzhHR9098jHDIDZAwOiRjo5Qh
d8qNFwliFQDOEBS1bwz4jB+/uQfuMm0hOLRZyObtShDMTA6GogZMHn/HlOWVNw4DerShMmjXMyLD
V3z6jgZoBT0oeg6EwcruYL/51OtdPXNuVxA03kI2n9Rt8iN+WAICl7zGPFyJsicGO79RC2vaiYqy
+eMS0VyEoVnTvmjqRzN+bOum8sbaxBIpkfEX7Xv+pcmQyc02Fr5UTKml934uRdeDcuPTzbnke5ZZ
swVVcG3Vzn0Y7792Sp37hgAYMza4RcLMVeP/U8L22TKvWk3TKVekeIkENaJpvW5O0uQ1XjOkP2Iw
fNjNVWsblZ0zWPYUmvpyrf01ot1n81i8Q0RItZHcaT5zA6MOVyrSqwUGHOQ9X5SOchTEnusPZXkZ
hGBhhUyz2Psdxy2pGZh58vDm/iPRaJRQKZyLgdz3jhPDPoyHelpDoLm1YUuycsiWpyVCwUCmzyIs
q0dtqbfPfYXZKPocK+dpuuVPQ1LUIfQ0IKW0vJ2rBOiNIh98RIFbf4q2swIt9ZL+7qZH1ugJDcu4
pVNsXFlwsuR9ozOMBKwoZ5xMUN67lvWC9RAC3uOcQmlj2cgTjUy5ygiaOD4o9NHNbaOS0z7BYx5b
yBfL7BRdhTLXjO2amK2/XhMppVFsCYZlTg/u1ymDI0UM6yKac/uUItXWkbXjq4m92KRM4jTungWH
fgevvYZuu1TuIq5P8liZg2okAW2b/J79DXudY4QjrmtMObj6QwwyvbQwzZZu2/fI6DzSuWLQ3nWD
hpHs4JLkiB06qdp4dMTfeoCrDIuwZWizHZZwP4OHGj56ogHRg7xh2IugYOgi+v/V9TTayCD6m+Ch
tmfahSxpJQFpakMTRqtByMW28I5QwJ3kfWA14q3tJlCBTQVXH7b3+K5ERCYqjb71Em/pvBjCzXDM
BKXtuZ9srObeLWscL7aPz+TYe1PHw6MlGmB5BAfREQShbTNIS92a7i0EtrQd8f/RCTTF6rLVBbxC
Rkr07ErZy9wYXotzSAAjQx7N9LcDH/8/zr3lJApm5Q69rjvlM29tqbByMaNq/haaNJGz4EPgIPRn
FUaYmjli67r0L2hwhreQEqGEenhAS9RGDNawsOmkWpwwqNHs97H10QNxcIybYF8zmgAUUmnyuh/3
ogaF9AlOdWPYk2fBRgAUixRLC4grWyTAhUdVZg+ZoLxLHdIPzbh04ElbFiXOXY5KNeLXg0RwacWf
2ult+e+jUTyRAbjaT3q7HI/VvBEZKc+cKjah/anJ9bx3QYEeKh1MIgTyQmfxfvClkE0/mOm3cHeo
30zNeo595waH5DR9F0kvsqs6xcHfD2s03xgMBrovwtI+VgR7slQgLovDPWzbjriNQDkSMQsYaN7p
/K/2hxKwLrfVK1COuhtGdMw11gPF2Zo9WmptFtfEXGJeQgKAHCu+tNFY4wGfbysMbExBKG3kN4xf
dCqkhHESbnAYcMNW88j63Ue+k+3PTy5u0axePsfpZBZnpfo4G4fzlBtFmZr1ERtBcfi/TNRu+bk5
ZwvPGpQb8vYdQV3mXOPknY0aD5E0dPkTe6mse67HoGfMPIKhwt9AdRVob1S9Dibl+BJ0jtUABGnZ
BaTJp6zRfZRsSN4fkEpvMWdYcXQDWRbhsXGGjLXHvV391evukeucFy7/KRGcT3X5GvxvZ+ew7J0V
mXfVDCL65yk7xV45IafSrWy0DbWp+VGQgN2WNfLwdbma828HoJ/PZrEEiiymRKrxK2KR6wc00ngw
APP10qsQ8xFg9s/dJ8wygmZRTb66jOAmKJyefmrglI5O7UJnFLTh9HoSst+Z1A2pwH8d4Q1hIaeK
AmejJ+4GQgSSmAqIn7hhpHMjbCmGQJdivIN2QzKo+BGZj0jimodVrmyDgYywA8WlzZCFoG7BPH26
XpSBlqpi+sNSXtM7dsxwTNHbjzSdOBygJVq1EaSyNaPQndXHpeG9eDl+rOsDu6F1up6ZzFI9viFl
+8oSOz5yQxzY4j8XZeIv+xnuc06D5PZQDObTTJc+Sp92juSMayPcbSanvsQ50DGa/ZlVukwPXlgw
513aTXMgPj4THAZtdWrCVnCxB/LeSMclLL/YFOjhW5KRjUIJO7hBc9RQV8vm6HFPtY9rQSQ5AxET
QR28G/g/thpFYSfRRG/44NRQF+k+/r8xMZFRpb+8In8ZC21jbMmkB0+1eFCKqLi3fSu/BM59Whzw
+SeCAMIiS0yvWcdluEDmdDuPE9bPRedfOr9thCe+njr5G5u4Xy+ChvGqYEmtquyOmk8Kc9ei6XYP
3yWvnKtOS1PWhO4QHP9saJxk4kGOE5s6WBs/el9obGj5+a15nPdegn8hRu9R1wPcL4ie9aU9ngUI
I4uY9uCd6j1guObusp0h7a4vACUQUvKdDczrTQVmFyvwXKq55GJeIWqMoy8ZDHoye9xdWf9osmJe
1aRLd77tofv0znAigvK4XMbfr7ZkLZtuOscBVBMCrR65DuTMYs7RY6Aikxo/YMr82D/uRJrxijj6
fSaOOyA5/2ZkN7eVzd0Dj/oX+dDTpoullUYofqMscrX9AhoFZI6VfHe9P4Q83E27z2Hu9BH9IqNS
e6uz7c/OPZCkCERmUJXjlPZQ9HYaecq+zK6lQJvYMmfIAT3wV4pBhTu/w0PVMgqMZge0a0moAQye
Po3TTnmGhJUuYPP7kVICMncRVvbuk2J5SFsvKtkyk7vqiZ677wo3NmnH1789pmzHrnBjT7B1ZqT1
lyjy2JKf2DfwoTHIfu6GRHCTCSVHZU3bQcoLm1DKCrStEVlbgDP3S9ynabhSuyx9U11Z1SW07SFo
/zvcXkKCeFGg7ccw1ALJ3r74mGTWJC0RsNLziW2Sat4XE5eivK8v0uGP5FCQVPYPx4RHCuJCRoAs
hRzJmjF9YV2eHxaWXOOhJ4wzMPOHeXp29SjVg8Jrh2gL5mwNk0cIVU1OZYHJySIGvFMxhuCuPNbB
ZC3GHFFCN2eaUgyVkoVxOkua90P0zTeeQ6QAqET9gHEXB6+6/WPlTKsP2yh+j7gMSj6QIKhodsl8
vl+KTi1lQlrfS/1Irv1gE22YanugRSZlo3c6sUQebAzrdQT1iI4vkX71dfoM5U3VEYKaAn9paF2+
+gp+gbhTZNA/ycZje/hcSGuGHQjaDUlw4bZHT8jRybZeL8NK2jwj6FiUcqnm/GDcLHakxZOSDTg3
FVBfx1WNgae8xefTIFUeKg5Y+J7BRGlB6URj6f8NxGTuXco+1hBRAb8V0MAGBHqOyoAGWZE8s4f+
484Qd+rRZhlUU+7Xu2IlmQDIgzdKEtSBfV5KNDkNGYvIjQfpQCQLPBviqWAcAwnK+r6UZuTNwHfY
J9VtP3Gfb9V3Uv2M8wimr/aHfDysRjiOuN4zC3K799oATyse6LPnpzj3/vxRZlbla8fc3LNoVV4N
WoWJSwWbltwQoDrnbSoQRPXAuPXAIIPer1GyOWcu4wJmgyPbhQachxUAHbYS4c7wTjflZCXGC2jr
oI1VJfv10q8Am+3Nodl/Io48eo0h0yBWDqeP8ivVP1B7S7rdTzQcNUbrbRdULLRZcToeLp9tqW5h
QhFXRPHokSfIsHUZhv13/gAMU9jb0J4vxpUqrk9pIr0/GSH+XJC0FrZfiI+gcJntNGiiVi7PWtE6
quNpnnCXKAs4d47y/IjMXv+PEFszG8f85sarWFy2U6ZyktnUyK8yPv+sOxtlJCHpgxrPy3mWLn3P
facoLd0/fFbCKbpOBbvYCzhSM8rMOrEGMJ6G9OetGqb3Uxgn8gtMF/F+6vKlkS+iuOHlZnoWRAhk
vce+DxGLVYcSYlhbbc/rm/B2xyh5cK1O/GYyh+8mrNIWOIxTxevA5iyC4UZBgOTBYrMKOG50sO8T
qQ728GZX2JY+HUmaFUvHLBggiFrqL29xJ1G7PoVB77HIUmHqUBq+b33KYJGahTcR+cWgyJfiOLS9
8L4butRGV3vyprwthXK5hEDh72DThp/qd23Un6rZzL2sf/nLB6FMAtQg9pEb9dY8D2mYBX69tEU5
vUVVw4VqfaO5f9SqfEkGPeBwNaZsCHnLzIw7+lA4QQE8Fe/Rv78EiBzAGx8zpqPMYCCegt47j0uV
f1i91EI51cDLBZxfCGg8KPwd+5BT2k/Lt9BJRKkfR+oMGi1cdO6wcHs0sA/moOC4m8mLF6MxoCX1
VBiom8aKH5MtnJ3RkGys4Q3Uc7kLPHEChUitza2gB3LHOlhGJJ/xlFUFSslKj03VgGWi5+f23JvQ
vKWSAUmT1cxvfx6KIJQuUyZZEPGBg78fvtviESM29HKVAgz0jpRRkN/WJupIcJ/eKvES1sfVtNE3
/jo2io3JtD0ZBMzbJy9wFxAtCObeib5sGFbPf4UeN7VSjV0pvmhJn7bOrFyqBaAbnJmqyjLk3Hqk
UasZtsUiUAJjFLdzelhnClfBiqF1Y8TjwXZQ9CRkG+HcyRdg8NXZmn/Jdyd2BC/UYQJ7M5Bs4/NK
zzFY2d4fcP0oxIFhYJLOvke5dms6ND4A194eBDWXXQ6oleBRejnKntgSJ8XRnBHbihq5UifLGlKy
eM/+3xiiYGFZxeKpu26VBJ58WjvqXtRsMwgX57fU41g7WCc00Bn/LM9+QYy7aobu5EIsIFMgq56i
KbxUrvqr/fPoDVs6PS3xG6quamb8km8u0tsEuMbz3WYR77XBBjdRVVDZ9Wj+Ex/FLK8ewCr0XV6S
MTZWVl43tYdN3hQAWoDnQNKkN1jvGLG/Vn+4tUlxaUQbzs30zuzNtweesZBXz60uyUbRvP/RGINi
pD0889Gb57GCtfRFlVoD+Wg3YEdXa2hWLkxzOB8IlnYaEOsLISKVv1c5f35/0/oBV9pP7xHUvtEg
Uass8v7nkLQJw5p4N11fR38CXrF5mqSGhcYvXQmS3oazBvTV+ZoFab3pkswlpNQHpdNF+/nmgtjX
TNEKz6orZhsfvXclccN4q6Fls6N9J1zfWu2FyCLdEoHbcc1vfv3k6mt9Z9PIOp++M1BDCr2F320J
FqLKmtFmk4A4NqXbrp/GIMgApMYrznL8vZ6pPgdyY/tlwmYih/kqL9jfvv6cFL2OWsWyQ6zgM+9M
EY/78MPvzWyy8U3xXulcP8dO1aeWc68oxeSJFxgHYNmPZxvxwM9e/S3AMageEysHRCXWGrRpVW71
qiK9fNC7AV3pkmT5CdmHY0eKXWd33Zx4rptd6Ab6N083VlwEbIxtnHBDbF1imNKfkWx1PLlvuKo0
R8PMikmw4kUnHWxvJiJNG2l8It0UPXb5FW3W7QePbhMBbecihk/aNITT7im/49CMIkVLXVR5wmC5
2aLKji02ZY6RmfrKtwZN2p80tLIecUQOjd4/KKUxQrCWpTw8zd42Mn0KGlUUKKDjfnbkmxtGFHFf
ysfVrfSLuQfpnHgzMANthXHTVe7R6Od1vZuDY5c2Dt0+PLGfB8hFi47Jy5MrNf/hPQ5B1e86ll19
Vo5hp19QePvmqjt/Jfpt0m6ZcTmfr7ahw+jUQqZbXcAKnsOuvIPw+dgu1HV8ZvaBLHjPqGHHOr/D
VZUp0mwE3dlcGvqYv/JyyWN8qEwY6XxPwzvVZDbahvEIPp7xkFECrcXSq8KRD119EpB3oa/C/7tk
L8egL3LDy5HYOJMejWyHF0BhN3zGqwDd22afM+gAcIbfBLdpsR79/onmFRislj+7eUlZoPLED2Zz
eE44X/kvg/fnkhavObJd+p0xVSgBBp82H2puwciUZE65OACV5WltdLwNILjwSe/LUWBEU2OGMrnn
nxrlIUF5g2J6FNm9eGfeKKhMaxFMLGTvw9Vhlp2ZyDP6/jQwvhjYDbUILMf+lQhs8c3/lVbrOgfj
pTZk/X0CZ/pe8AUzsHfkDYtqaJiQbvDCrUGvlmi56T1bdwD0rfBunf3gef5PPV2uf6uSNuDwmNQg
QDeNhTwS9L6W0TGpxxGuQveaL7DBg9vNb7lzLLbVVIkONKGvQoiR4ha3FcXHQ9DUqOliPDOATM2+
msjtV5VrH1RTXjZ3qfacCN4S2cwYuZluZg7KD/dRj2VEwNKmLAmEKK9rfd2nZUgG0gU95V95/PLB
wWDQcMpu2x+jcfc2fKhyytmq3N5dgRlLzmcDm1Kxu7zwwqnPtBh7jZ8ZFkc7hkdISbZ3DC8YrtQv
en9QEH8GJxNDHOkS6WOepDPzvpHUaK/qtqFNNOOIXFUrDebuziS4fNDqKSGub9ycnKZywB9MxWdw
oHbO9MK9cbya5ghwMj58Yzip7j8DccFYQE3E6ZVNVHRWcIQTzZ6p2XIsVHOZVjlDRQVGcGEJlWh1
x6rpeet6CCdO419x/KFMWLPtrVR138xYEcms5qw/t4fXxLeZh8vQsmrxCATkEDpmGpo6DqUYmMDs
nqWQpD9SzJM2t1g2S/3O3nYN25Sy4gR1/7qt/SCcWiYqGJAuSsHPfIMpr700FOnCudB5zxvhSn8m
xFCmvzMWcRNvnnJ0ZRCSa/2q4wBXs8jQfzbNPPPOj89ZFmqKBGXbCDIKW8cw5FmU8UyfMeslsv+H
YOsEBXGyl3x612OJ+RjjsnKYQ/t1FsOpVQ869c1h2yM6l+OcMsATg+FbCnhGGHrK4Uz4coj4o7uq
JAh1DIxgU4ZpqVlptf2MoJocxOaK/1ik1N+3lJ5b5gPYmJ5CsFi3Ebzlq87r7O+W2UBu6w8NlyXj
lBwya44bxfT0qPMgKvxvYaZIRxR7JUpzfXy19UTx0JHsaA/FLMtwqsaITk6gUZ1OAjMY0PpQfXr2
dcYfDdkz2vws40x0WFBbhljPksNzFI+vEqBxWSDbwKXyupCcwUssmsO8DXSMpWHnSSDHjIKJKgJO
e0DGhZhDK+h3IRua4zBmNtAJr6O94eW8TSqbpYFfPBJwwn8urmCQ2+g7KxvESdpw1E/cqChbS06F
KTgn8zdlvUdNo3TxLclsKw8C4aHJwqKnhiZDtRA3ViggHOGauDsuO+T9ppAm+ordnNNoN/tWLOC/
LJaQrN+GRoSkpM1r2m3qldIw9qLebRR7bFdWOpXiveAUa8JbNuSjzswwzBRROWXYx/qfOe4CkVtz
1ae+osIuChC//Mrv1zeLY9rXZKIzU+AKxegXPQ1sH8eJyjV4RIHF4nv3vZfqfCXbQQaK5SdGjHh7
ygKlDqstqq7jqFrvFeEZopFczzFZ5ZXKwomlDQXOXetRhSSQ7psmS67rGiEy9UwdHgmHjAdvSRqR
mJk/6obuRmo7em6gaMBwvqNMLhjle52MIQoB7MsHoYPS3Z+7J5c2nqel5EAsMpYRd0GIpN1yOtn6
sLYeuKZTUEHQ4QoqhzgFip+sgGrZq8vpsRgOVdaueFE8FdW+J368+5fJzePTGodzIfGUMgjDU711
hg5Mper7cLrpPGF/9yGbhrPdDI0bHjWEacxnvj2uuWHt6YjpeO4GhdgvM7v+nbHFOQTDj59Ht3OL
GWrrNack+sME/LXMXuO7w9jsVGYSPvcaryhR5wXN05vcFDEgSR+BZKf/4TcG5BHLVAyA/OUzy1IU
68c1OpzfNjMOwKz+T6tft+Kv9DRb7pJzAYPcfviDggcjUPpJnUqyy2zpLEM5IZF6dBucLpfvI6wJ
q80CRhPcb+aNGK/ItGCVT6lEBEtxK59LUYOoep1EnYt6X2s8WVrJMMSC1UFgG6w5iL4QWLojXdFq
1n3bSz9skcvaUiJAQqfvP8mdt/C6wcWmeMSzE8oaNSkFxWh1I7w3h6ThODmCXnX3zRdRMcx/tSb7
ctaVFT05FbVFxRH9NMCOdO7UAr3UGBqQuDWLC9YoOMSrGdz7HbPX87kGglVXIXNU8clq8moyLMvA
m3BAZ7OJPIxZyvLAnindMOs6/qjoIaxWQXDJqFKBwmcMgOiw8uCi9JUpvSVsU0Oy38kVvD+t8RCt
ExtagOpKozdvs63JM8lH3FmXpwLcNi1TwXPRb9ka2642t4JnKuhCJv/HYn1UfNhTqNMFNa0yLwJz
cXwAa3sDOTG8hGWdhVqr7HgTEN9gnXuFIhokmm7wwQGuEsc13Vun3vK0n4FUMafW4YvjTsch+H7N
GjJCCR4+LR2zb/9h4uw4+ehRUgIGuotkzenbpVTj8Ev/vxpLYV4aEU7VvkW8w3zQANMrP+t3pm/Y
1eMv6LNf3wF2GkJPoEb7TlV9eOlpQknWJamPONz0CCTf47C5c10maDF+3TAP/XiXWnfszPqMZ0b9
rB6NZsWGA670de+WumOAzxyACRc94TLsZjtSSMJibVG1XuBoh5e9kMTq3VhE7eswyzJ7fc871e60
6phhBgbrM+pYhJzpEhHH/DXGY34O6tgdHw43PQkmNcq15BZP7xZom5BX5964gOk56j0pDWus9o9G
+2ksAmQVpWRWT5bsYSJuNLXwm3o0iTzn5T1+0WW+epmi0TKhlecxmMDAnlDz0nBJEreyG+/s7bEN
4GZ8IGh6+b+mNUuOHciXSAnYxE/u47om/AXE4l2kw09BFCmuSJYYEyyYbgFFb1ZYEvyIoHzL448e
dguKSdk9cFet2885hk8OkrhlJNZ5tHk1GCFb8UV4RZ9GfWMP87YrvmbmZycxCDPVUV8+eMYz1uRp
LWal08VNeq8eqb/Ve2O5UuBWXfUVjeULhmh4zVZGqr+WMf+ZQ7s7VLQqcJeeH9luwhDnwlVgH5Nm
Tn35LGh2T963lQ2FyNTpcpmISBzOrduNlfNn3CYMSSQeuj5X4W9k6K7mf6HX05gVxyJxPjCJFYyA
dFxRRXutdfDKNwCYLTgWPRMyVqyCdAMWzl59YfDWdV8v9K2Z785ZuHksvSefozUKp3yXTpauytG5
63lj3JXuBVtzCcTD25UHn4Bi+70uFfdufwrbBjiwSnYDbqwm8X5EoEhCyFkDK7ElYlHCwSWV6wN6
eVBfvJpc4EwOMMcqUyxw/0g/e+qWRrh99nTJ7UZlIHbPAavx0YrXFDM0G9AOAVAEAMjUHh7cJtU3
orFPlsKh1eQC/kiTcvNpGeGDHB89fDexuFF3dwS2H8qg0vHLj6/6u4zn/ROWZJb/nBPcrspht6jv
lJ6O1VHrFq0CHkKKoglnZpM2K4R3gNeeoV/wb0OJ8tmUNE/r2S/969lkdY0Z9oqGcOvOrd/K4QMn
nfzVs0l93OiQFMkkjFYuDg4RSud6MEVRWlvQbVtB+ey1SPpjiipBa0BQCbzv4obopy0PbKs0n4hk
dh+G3fdmHLk0QBwhaFfv4zdgDJayV4E8mu/sypcL1vymleJpw70bsF0Dpmw81/3MB3pOHttNmpcY
RX++ABYe/52upbKMQ3+nQnHN6m6g+dTco5YfZmKx+aryE2ECggoiRc8T5ItnlmrO1iMmBYxx9FNo
PsPkIO17aB0i1Lo/X2o7eM+y+SsKhNs3wDhuOkjuabtYkYBYRhhwrJUUzkPFhDqsvQX7Cd19+2Pq
EakD3Qx8ak+aBsOc+vf1nrVwbUwEPUJiTw2sekU6V1MxQFiYi2XqQQMLfeD5vOTvUXWzzjRF4qLE
f3fF9SmgYe3AKQw2lZNo3mEfNzs5wZZs6QU/h6oGtx8hT4ut0kb+tQYRyhLHm84t8QpqEmcnYJ5V
rKS7bjP/EHH3sVn3LHdEEPtvXPwEzDq8LZmepZXCd/nVigUGE1RztuDubQKN6rrS3OJrpLScVl9F
d6C1gvAPxC0QTDhVzthIyuO9uLQSk0MVtR1nQSAauR29tvF3NsjzpV+MaEICjrrx80XU/uP0f5GG
hbEGEpkXz7Q8pSWef1xaLyIBIG8nBE8RBytsBmOeTAUCSZOAr/DjFwCD2sfs/4h5Qg+ibB8hEFjv
56EU1gou8Cb5U3p+/AhUZ+hCIJW/615gP6/8VKrbihp7Xaf/ARFz4jZpE+/cUbt+lFOADOQBr3jn
+prumSkx3ZTn52sDBPqh6j/Brwxzem7d37fN8M4MLuDRlng171XPUqBsi28lGQpml4C801KL+8qH
y4/vyP3auz4b++X9MOlkCcDmzp8FXRWFbZltI2S8QAZjcZJwZuCDnnY8A/kzKD8xch/Pbuy9NnAv
apXf4q53xbQ2/bFHYAw0aDX2+ZO18NHtTgwT85h9yuhSB+hjtkulICqLlX6SHFp5ttnXJESPbHPj
3T8rVVGGgLkiQZgGvK4+mbFxd6DRTyP0KJqGCVUMJ9EdxbszzEwA9XsH3eYOmIrZep+xbWKFrqKl
KRLp+EAkASae9S0qckyjKBy28c2S9gznUWt+E07Aqg9LQuL9C0qaj78Hymc4gm5JB5Ra0CY6mUJK
QToe8uov4unga0b89H0TRZc5ckix57yxAJp6oRQ34SdIwJWrOjsbhwbyx30PGemiXP53AgLc1Cms
AEWDVWCZyrNg7Wg13rxNk9z+Y0glXSCGCSyiupON8HdoHHF5plMdLQ7M7BY7PWzEJ8XfEyv36hK9
NXgeBFysV0ykbx2WeO/RKPeG/uuktZ3JbLypo1nuDHQ7IQyqDoxa++gK7gzbP0F94mS2dsieNRqZ
/P5EJ3V+T84wgwHeI9hEqVX6VpVYT7EvMiQjYFQNKCGSbX4vOzbgu6ocX3ZjlXooCqusGvKkVPBT
Ny+40vNkZMLrjE9yaV00DMFB0weYxbgha7q01qLvgr6wmlUB/nvAB+Cb0Mf1O9npJl9R7xgE00K3
Cqe942JktGLDxboPBBprrcUx0uhCIlaoMsV56Pa9M4/ABNu2rRrYnwu5n99Uyc5pkLn6kHEEGXBE
7gCD5vDlaQDwJcFaKrp/qDolxtsYxnTGyWGgB5M16O5vbVNWwchnTAccmxSi/fmxP99LAoojdU6Y
VwLB+uP89AIyIpt+Yfeea66NKACX5gB3fynCs1klGMNUnQqDXS6dxZUcqRNHnAwa7nJ7L8ftXoUM
mfQuM+A2UeW5OZPAHYnHTXbSybjqJqhGLkeilAH8z6CAL90XP0loilZ/JSKavdc0lRMTtqjQ71+r
HoVtTYNNXA0XMt0G0iWBVi1gsgyjTjVIcK0g5PB3q45B28VPx9uCU7bRlKxyPlt1zhmMc0akMZqM
0EMM2iEs3ylt9T60HmcspJ2sNonu/fo5GVKO8WRQNmK6LpsXrA7Iib1XjeJsW2hK0MYtsBtWFGu9
sp3iDIqBJFqcJF/3tEI9b/IhsDqnnXcSecEbyznaJ7RDODJqmOlkX+bXLQiFWpC2iEQaGiPmeugA
6Qu275wa3cxtr2Q8FZYaBUV+gsE9wGpNT2r0l+ovG3CgcxUsgCS6uSzNIiM9/d3imJS2MaAsQ04n
9E+mwQiJzvWk04TXLhluEammrKsPz1Z/8UUU+/LdPjbOPa1ku4fXSMM2PC+fCo9ZHmQ/gu3nXXWO
DybjgXEmDkk5pGYCGikqq2XllAGHjlvZR9qSVRjeptKco1VPjpCQzZjBTi4gdqDQK8K49U0dzacd
c8gq4VbyNXmPcLs720UcOfRc19ACO9L1Yb+M4uuAKok4VjgghluAmGKG3/KApTwIAwPJW9VgQ7hx
mwSdXjcyIf5Qhicqm/xYvnu0/b2D2IssXeAsvTvgg+Fs88/2ZfMoRjG/nDCBudnFTHDvx/6GTg9I
9sYXKyA4WvlqcUBelFXBMB3gDQ1wtQnms+/Md/2R9t2QgclDol3AjizKFh6vdZd6lwFHw6a+u7VO
6lkTMZIooKI822w/sFWRj0PI3IWoFFX2p/+u3DNb68At+KDhOhX8TjzZqEZc0zcl/sr1i/bpW6S3
ubwVuy5N/QGyUnedWjILxxkOGwM79nCOdAUhykbeyKeMVMIzINncggTHzflVpqA2GBt1wtatesp0
niPdX+GudN8txMogv4RxarFU7mA/Xd/rN+OL2Ik4FGUAtnPnoYncBTIksexiqzFmPSi7Pb6K4oTg
i2nsEUVlko6BdaOw09EOmO5hLlfRsZbrYD4ZGH37oZKajYzxSXP1uPjmwr/JvG6lMuYM5k6tXkYH
WeuJTFs7/Pbz9UrbojJUCWFpYk38vNrFbUZgYGStuPWqL8ZQOt5CyqXXyIaHvuq/nyed4azoSRBY
4i2p2fRTxSmN4o1wQvbt4z5PRom604rOMRV+2NDEV1RZ+1iWLyo+xVL4IQM1AhCS2vt0hiFvOR2Q
9q5AzKo+tKj0Z4X8PUc2m0+S/byKxRfceJyBxh+Y7hHt3/TzdGQzxN2vgTRm3F3A3popdrZ7rsFY
f/YWPGhaGlr6b30Wab1HqP+KRjOpiPowL784b3+tE/MfCtnN01yl9ayHJ5Wnc+aHzX5pWpc5v4FH
mzi8VrC1fywXHxsRBP7W+6lnmIjpvZ2riYmfTaccr+EW/LY6+IPsgUhm2g681PknN1gA1fRCb6fn
XVYrHOz5/vcIKgM9P+WfWaDvAreRwnuVL+NgmN00qWj6tNi+9hLCDqUjpOMGaTCRA3mok/IwqnyM
hOCyH7e+EKis9VluC0qzak2J+vNFmtFsJcMRb0kU3cqHcJ6KR5Z5M3EDvs4Wl5fCskHrYPJu8RAZ
VFGovgJWiRde8wxLroUGTEA6i1XGSnzAnRYfkNeoe7lfMZdZsNjQhiv1m4noo9OOSU3nL+3Ens54
wrBPn8KDB2eX7Y1rF+CPC0xim1rQvsDh6mYJKyNLfdkEGE/l5Xf6DjZhSmSWOCK5JmFX4AXP6yq8
QfpducsKHuSMdRojIM8MXJ9O6bNHFaZjhYASCqRlsKKcEmANkjORvuQh+T0S7vVMZzDksdPYhlko
xs1g1qeDSnppl4uIeAfHqogYJtCgUhMG2NkBwCnaZxqg0i1eLjr8thVu1cjDmaxrHLCoxpTgPjKU
Xw6v/KNyW5gZVLklJrpn6ubAvFSZ4+BFyeoONwZ8CySvYBOg29JJUxS1AtdRzF7AEwyYJ03p5Vhn
ExXfZ+MqnPrvvTmtUGFmlN+EqRehLzeQXvVTEC8m2/XFzITdF7eOAatQKmfSYmmKcAaboM4ZkamC
h760SXB07lIbwkFvFp1tLOMhoy0tluqWygpRKCerVxjnEG8tlyyKADXPDgT4NxVOmLI25mYm4PwL
lDfGN9iE7aNB7c20l22Z6rWFn9RBeDa9ErnBVpx5C3Io40pmiKffI4K+QPdUzBpBKnUPUoHWTgHp
845olwSBAYFBeREl67B3hkloG9dn5YpNYqXLFeoVPiPe0ZTvXCiF4G0sHuDfrbTrJSRhNTgusc5Y
v93kkUK+CV+sDDnNN2YIAgaW5lg8KlhLhWXcMwO2JGJH5twvPm/IaAlQszpuQnZ2jpRleD5crKsi
K4XsIrj6BMW7Gfv8J3A9QMLhwG0t5JBdrASB5PKAuhdnemwpGzcIooBnqMI7X0GHsPyPpFJH4fjs
IcrYI28sscG3WKWCkuUaoS6o/MwzZzVKFtUqwbkmv0qob7NomRk8a57Kx3NnJhtNKDVySeUrqTcR
Ul9f7CEzo73/X0/vM7XZospZDIXJmkSOHYcIidaMLtnuU2+jGIBjc4uCC80nAL/JRt6QBfHXVm3G
E4nk1cNmbHA1qWBE+M2SZup+xz+Td1N/cF4HTGsd2PS1Uu8y4gAFmguIlpavNBvMGJn0WThLHOrz
5qFEaQuqydsIUa8HMSn0SW6fv0jmu0kNFqavKvccqUCI2YArxSnnA+63KihWGc81ESuOkNAoVeSu
Hs7/K8CNIzqPioX+8ws6o5hi6fb5KErwvrUpa090I1J4sZk3v/b4j+cjyWv3qBQ/CMnSJ2l4uPjX
cw8xLDbyzJCZ2214zppe3GGqZj2dEB5XR6arcM4e+5jm0e/tdSJ0VJyUK29qL2FpJZ5eulTig7WA
OT0u0SJv/12FooIvBWNZtYCftKkeVfFW/FWmi11ga1tH7/XhgwjehqXh2aNzDIkp564Fo0IkrtiC
n+NQUYXcL01jKjPGCPPiX1+1i1o4NdAnkb8vzWuJpqlLkeKYsugCOKHLzVuUiW8n/Po5aDJLszLk
F7XWYEEv0N9sfON4xfrFdvLzK0c2eXpbPaxeDSG5dzwf5PBRfeMBn8ujoRnPfxJEylCw3jmWEQUa
Sstvdj6lYEjwVV/X3PK/kwEA3dqnH0wOVjHQRoAjUcqHECQaxjkDmBrSc10n2hQ0bgPmlawhMba8
sZUAmcEv4t54+S65bngH2YykqUUoo5F9lRSIvUvi6wv0XxlMoHN5TqCPmEOXieEQ944fujJzMl//
i/wSKC/IrSDmJsZi+KjqvYZWbwzL2ptwiueingYC0GCRC9o40tGdE8Tup8tODpDcoDH8BRB04qXX
PzRvOO5o5qoA+Nnu7E0nS/RnDy0S7tCcQXTYWrbXCEevhVtKzJXobAzxI9ffrWXLJGTQXV7tDjz9
aAP8E9gARbJFg5opGqMlY9MU/pp977I79ISDHSYTujvFl0aUZRs9FOQG05KR4AfxkTijpXGCacpM
C1Ikytmem60eCtbUfkvn6w9KBMsQXZkESDNsnjr1ptOvu1i8fq4cWCaIquFYBUy5AwqLuZVTtERP
hq0BSMc83nSj/OLDF/CHLzjbid+0Ex9DEgG5PtKcjp0CTG9gz1JOGQx6rwyj4hB5sl6VBjra7oil
h0ng1HpubkAATiQ+EI9p676HKKhuPj2wYgkQWToCvCsg0l0H47wmrN/x65yTWKNEMJo9aBOdHUCE
DD7DeJWOl2r2xEe5B39y/rSJl6kZUBCM8FhprdOTjqRrje/d6jZsKZihRL1ZpcCs/iSXAOz+YtVd
Nb2cX+HiJHvnBP5J8GwS4dAs69hCjt9tdEtF+KsZPKwwUw7klnOmLl98fPPo2cq9mBDzz/YY2nOv
+U1q29cCWmZltNxXmUej8kQLyV7QBoBg0j3FM63mxLPiWWJuyJBRlv1wtR8cqBO4OSvpw2WBie3t
Rujtg3683mFzJG6qgstYOMGSbYf5uwnc+HcqVv02FtXowcngbyxg4KDRM5i11q1wUdtOqVB5yTUB
o15axnJNvc4RHnL0zFp5LHrn4TYtZ4EIMHk2j9H9svUr4uwqfpXVdycSJCNjVbGbISIQhH+miIvX
XDVMqGmrfDmRdNB3udoBClUMRL5AWoALQaLcxiS800OBcPHWit/mtMpO/Uf3c8guiJoTksWKhYri
zCCMsAyEahFjpoAehtdwkV5k4bAT1wk5Q5GVQcOF7XhE3Zu2hWcIj3uC5L7yGBpByZlTfPHeR75/
2UvMnqh0vYDmFGt4J8h1NULpBPHt9HgU92P3TQUCCwGIV5gsoErzofXKJVJZrNpUj6RBWEbaaux6
u02dmqIzpMeQhATur+EuGpQEtC1jc/5JI9JtKY5VA74CyfvkJMuVqPyumik/ZhrV+9jYOV2Ofo8m
pgYreztuuKgW82rlRjK62Hv0jtbr34sMLdp694cxX45y6jNBvoT/qLAMOKUFM1TqCg0X17r8cniT
3IYj1k6YQC5LfLoiNH/sj+6Qry7quJbvuQH0+5jjLPwDvHjCBtNw9zejF9/0kpeXNbn7f+FwhyuL
Eh6+peqgYd+XyTzB+x2fM4QgLt5gxgjTskwMTy/jDEn6h5gb/mOBzoodJU5v9lsDN6PjAJ0QobeB
ZSG/JJfVM+XmuRcJYXNLCpKQjbAMxI8kpQJalYT1eWzhdhdLmtdOPxDoxgoy3ZdvQOpupH+qwfEu
vHtgQXKCfN+Mnx0mJMpOS9f1aD0CdXXvADNk2dcl7nWGU3wPPdxUgIXSophJfYJ+F7ePePgAdql1
phTdxFum+RT7NxNM45UQ5ItJjnEZ1LMflIKlhpp8ORhGmb2lw+gtMwcRjVS50h8MXkUf3L64ZBrN
hT0QkGPZ3QTCsZqHhuZ8IWp3f4JDpREaWlSqAtxiWnBNdLBKpbe/VCaU+mKWZ5Bm4xN1+qT7UYC2
hhwl3+wkfxSL9xMt/iwj0OXuErebxMlITL/aKlfaCbcDxjhKvyRrscLf7N6qtn1MoKowJUE71bTW
GSUxbX6FN8Gv4e8Cq7eWZUtKfxGcW+EzqZfBkZlMOLFApXBGPduOvaw78osOzyXJWOdbiq7DWigF
cmEJROP0V+G/uGnQ18armREbQHLCiIAbfu+VW8KP4Yh+IXSED5ir2yYGr0DX5gH/hi86Jiv5Cvd6
bWECOJQckRCrp+iEcQt9dKKKP2ffdUWQm7B2WKwiZnzSlK2bnKN0XDoxymbosHBP0KoO7NruUFeN
kImELAOcKxszMeNtQhHSyqmdHlUf1g9QRkBZRnFa+nAmz3nAVsB/kx4P1R01PRi+SCXQciibN/f+
t+BJj6zEH7FC8vbFMXKjTJm95+9an/Yh6lZSL0PFGROqZm4wp44pssRMnjzSVMvvnAjW1Rr/gtcP
ON2PDfWbD35BXXo+riz7QzYH7ZdBiiNao5BHphHns0LeM175gtXe6aGjBfSHN7XjYzdlcS3DBHla
4u0PkqYAXh/Y5k4OZRkQatHP1Xb4fw54rpm9UkT1LfSVJQ0c3NTf6F/HM3y+0Os9fg6ipUVmHls4
tK2jSZ07Mevrh+8RvDK7nk5nvYyoDfiPi0ExbuSRB1h8C33S97hqAaieoClbWw3Gd455Adm3qcGQ
B2D25Ah8Q2XhxMrLuzXsmHeBg7hiKYU7vvdY4IGUwdT1AGNbck4b+qB8DSLlt/rhptPQHHXDnxTi
3GLeZuBuXziBPLmV3jpbeZszCOIKb4SLctYrXK0JzMzYlati80wHICdOG4VzWO0kijFNPLbRgN/5
JMRixsgmw635lTq/6IlDu5AlNs1LZPqsnr9TzOuQFm+JjZiydbIVpvs2AsXZWdisnirMegE0LFK5
m9mvfYFKSKQOmTMaYimPioSBLcDCs7e89gDRs53Iznd9QbO0lnrnuewniNnrHm82qCgf8IpIkswI
hV39Fy+rIHj8a+ndCceW7wjVh5FYUwnVxpf3rsIbm1chA0uuL/+hacAWnqd8eQeQTXpUZoCN5usw
S78L+AhyCZPXM0Bxoi0UPbPj63/+2ZwxBIxxveb76pkDMu9wkwaKaL3VaNAivlR8N7Ydii5DooWB
j1tiS9hz05twJUPxb+SFRFTMU5hK6UqUE4v8ZFoezR3boS44bFIV8V6SQ8zmE71wqoZj2ZuqM92O
zJmE0CazfmQwIK+yWykKTZXxzPJuIjn1oghzlDUWL/8EiFo5w11aR0lcoACbfjjzA/0OIqt1s9lq
m/9rqUcEfovRxivuwGKb4dmSCj3gjJXnjXXtp+WYCn8XwmkZnCmPczynQyiQIg0gx9q6p/TsGmZj
LY0Wsg5K5tOOrZ30FhoAbmbHcm76d9yFYq38EHTgnCaVJtXUN9hh8RMbeN0Js4bpCRFsHuyG4Boz
Kuq9IxHPnC0FGv1mh12DFa++vznn3l8fkxd8U3qidCkEGbKTFD7hMGPIHg+s1ONR4NSY3DoN+Dcq
dQ8FYeIWqOMJStAqV47xWO5OZZpTA59KWNzhLjZ6kC8B1FSBQ5lYqhTTgPZFay7i5ANji8ymgmEw
ehLhGt/dx0TEKIYAR8ztUSSsyQNZ8OscEguMoI/Iqcw1/3MHK+0Z/IV5QN7KUuvPbKghOSno4qoX
Dblo02Cn4mYkuckoLSKsv8CLB5YGOqBv/SKpqp+8w59Xnv5BCmZ5aXz5nfxTtw6s+hRl9IfHvUhH
pHjXeurLJCiW4zx6pc4y3g/Tv3s4fmqgKI7DTO46UuHRbdmzoICrEVK3/JuxeFH0dL6qvK75InhX
Eii/exiCdlqKujeLdrD0RX6QKRbMOrUq6ajAYcBMtoG0zxLvuj6PxAgmyMyr9w1gDPZp3UGujj23
1OJaTijEWDaN1fREK7T0Zn1H6c+pZTnTAdywq2EBnKZ257zOlUPaNYuYRBjUtQYmkH/ky5Ci1Kqy
I5wuUWalH+11liPLHdYUUomb9bfRd93Kq/g3mQ6L6pCiR+Qotqp0t346rLjhcdozVI01ilwUWFIV
h0VlZEwAYK5cZkO65x7p9YqN28K15UtyzJ72lfZQWXC/qhpXZmYU/Jw4VoM85/0KFRHEXXysns36
KFlF/8QtLwWsGCHgwzgbmG+ZEdfhF5DREXATuZ+saUjzVXAPnYCNochoh5PS2sX8qGhtYNZEuCG2
H1TD1VCZzmzsYdb/ntQS3MaT7xgDOroXoDvC+Qd+23ryc+PIfX+EkP9iomKGiw0yapvtgN6dxEbw
UugJT2yMp2cgSdwHynMhnz9sfnXUw79uQm+Q8G+RUPmadjsTi23R1SFYGXP4zsnvOgqkVOe65qNH
psrxcMbP2/xoWw5cwzw/jrOGymN8sC/jigYaOeFBPb7SrXLBoOXQgiMQcD53zEnPDxO7dPSkopOP
lfsJtfZPXgnneciTcwCCf7SR6zqGRKP0ydkukEb5ekpQ/CnzIReKI9hAWjB+4/NclpHx94MGo+vN
mQAfq21klcoaiX33ajlZxM8FL3CzYY4rDS12arfU8qS3G7y0yB7KnDsgbqW3gNv076CmvSnjMrR3
Hkzw+0/gcjE75PLM80dl08+8pMafRpjjW1bO3omSph/WbbzLEYKyNQbKWlajeyd/HVdb8nrqhlxF
tjUNL7T9K/VAvyg1iq1JKXnQ7c4hyQrYBfYjI4mwOVKV/NphssI480cp6gvo5rfPH4K4Ym/oBaOR
+zvw2D8T8qIkS2caIBfv03OiQ/N5m6TnTX7/CuE0ZJlntiA6d16FruZrkamo0+TSov1KgTprvCSR
yY7kVTrTevuOxqka5uR1mnd8mHEZibjYP7bEpJNpf3z7uQrpafyI1DxuSQ9snQzLJyypQGu+kt9f
vkyf2S73JQ2cy48nkb5AybLl8pqHBbp98emSPMpwcW4Xd35zXGnqHWvdh67hhMeudoRbQ7lnVaJq
D0kMeaSz8Py4XCYebQonj72FEFN6cCKTev3X3us3H3/WGiBS2jyp2armA2S4ZdhQpkDFaW8qMgt1
ooIEzwo7svsEMuDyOjxY+TU4KHvcSu+LD4K4QO2gZEQc8Qay20lduow+zzzfh71yaYFIrbr3mmrS
cADtLAznRmtZeKS7l1UyKmkaWz/JbG6Jk3ddLEkhLuxHAKYPj0wEikStRtwTE5JttKFSuPJ2/75s
+Mwl8CEEOH7dySVbQZxrjxGhHLOXz5dixcir2J0RaV6sAHsGZMchib6leU4TC+7JOFnUeNKDV99U
xFKiNFJ28yqbqbhyYmESI/QkWl/M66018pawxZ040EoBUXi16PpQXd1gZfFznqfwa1SvyDwvqLTK
u+BvbWyC0U84eN/IyaBgNHB8jrCBBMjtCCYeBMdNuVPtzbQA6QL31Kg15xSVJU1ahqvPuaRRWNTY
oQk9gh6Y+J49J6i1J+D1xmugvGIB6DJ0Q7KxKlZwfrlI42lhK2y3b49KFzBRLKFmwWYp9m5BDu+l
BWO8i+B68wQoNY5Glfpjx3r4DF6jI0rqkFjc2LG1gfETnxrwiDuq8Hbowu1C0ZGdL38oZ5qHaRfu
kim5sKzckCQszoSFR09eKRbehL0IjVzEizYXAxBTtNJJRYgqr7Wvyqka3Ib/tW6YHg2bM95/cju4
gxTEdiUsaArCHpXpNS902mlH2xP3CiukzqwFLsv6OKJyQ/dywVg8Dxs/w/Vrbb6/n/OuQDBwhFFk
zOR1bV3leZ3yGlHABEe8WvVgU4O3inPTtLVXI87E6Pg9pgWB55ei3L4767Il+tmmT7nKrPFk02mn
wkWm6vFWL7kzj0Qsqb5tY4IpvGZxgJ0r+JwkFvg7V0+h0o/WiXxPqyzjqIC0sV6NfXFzQlPvMdLh
fwwFAjyU8vSzfXwkWlKaB0raJGX8ottCKTQDNMQkgh+3J1ztJELXaLZBRBMvMzxJbgtggiqhEzO6
NsqQXydeqQGW/eJ5vxSt/CeBXCgvbYhfPRDE+mKDa7DhPJ1ubgBp7IXB1E8/sBF1gyMrtDByFZa6
hIwojdtKEhokfmjZNxlZEqvZdH7uEhFOQOFfMP0X/6aPFcMqXu+Xu2tzDxDPMA7oeyrcuMzWwC3b
d5/6s+MFpEWbMvy+KZq43MdizyqvGjFPj4V0jyJHItHWoblD86dfbLbBPsjiHDF4YAO7CFZp4E7X
bMgHW4T7fLmO3CKba5wka/mAuro87VsIhF/ZlzwHaxJaVIpPC/UC7Q/c5fPxIb0aECg3r6dB0pia
5IRSiqpAtRphhQoOE5Yv6L1VCPWsVcVK7wpw+r2OQrSmVLIPoO+mnFyqXe8n66B7pdRAKoCtf3il
fNOikdaetao4990pTzG9ItUEOIwFUbsIZ5QQTDUivKDjg2OzJXawDBK4tEja3Xj4v1QtmHi/9Yds
Ndi7nEd5OcPJNFJfqKLDLjc5QKOds2O8gku3jw18vvM5FBAIZzBLZaLsCt6h29mcr/949xpL1bdp
vnFxu37Xc9cRIDiiR0ehmwGwE54q1uYWQUjsjU0sbZkRU+1dhgjYs6ekNHdvIfMt+Ook2TEVKRq0
fw3yovVq/UCcJ27pQJkN1gN0ZyIp7yp3wKfNb09aH0/o+DYedPa35EzTfGSnzI4IMTRhAwzhxVCU
wnyL8UXjVsx17Duea1JggifPLxi7HhmquJQYH/w4rLIFZXxeCpk1d9fDDgIU0J9cx9xH1yLRWEsZ
rANkBCn8nPruUq3FLUaZ/ixNpGNQktJANMWYbHf47uH4bRIb8dpdbp7ZwbK84cIT3vCAMgzx/Ub9
4+k2lqcbzr+WFEMtvRyHuiGuh48BEV3pv6kkdbqs8aSK4G8lJvjf+Sa8n4y6DtEfr4xtwxk2GuOE
8R7FUXc8auvTN0psNUSUmxg0xmYH/Fns3V3yz9oEhUT9onpIT0uGTtVd+gEP9kxWVIsd9WJ788Ij
xkuba7m2G/5/OEqvjv7StMsZz9Pogj/I47YzIYK7YdP9wmNEe3ofMDXYoxN9UyuX7RBX4Mud6IWg
NqNSQswsqDyFlLL5Q/De+LwPI79Bkw6JdQ80xWoGXyxxoMTRkKopKGqkWAYNMRoOdkWFLf5Gc7LV
Rj8n3KcVfkLFXonZGU0oRXLu5Y5LlzDSHBUiD/+woFYWrpKG0ObMKT9BzS60LB7sUdj61ntNLA+R
6kMBwTtXuhEqtI0hQybts4slBH5MUBtRTGLUadMwGwn/za3zSTrkaDxcU0DBYcJeZC1kIRNvO/jy
w63j9kOe/WPz5wj025Letq5EwOrRGpaPU68/gRxj4kLvZevxNi1rdyZWnlH/AqCqR1s5ZFwWm94D
PawHwwroz4vPrG5NXVqNoRT7q/JoW8U9DjX4qOpSEv8sgaUPeMpbTl8y8RwM7PyxyAIiLOuo0Iup
RHT8fNcq1AJuKJcaUj1Q0bubEtkXjWNiYiwSFcsIHn0Fe2mNixb13VMq71TvWytwxeheYGXzH2U2
S8dYLzbEyiI1d9jmbZ+3PZBAErWeF4LEw8eoceH9LTEQR1Ax5+sGD0lz3sVRskI+jzbuK3zGPIte
wJwtBNeDj3KN2dNOaRk0nml1vY3zzcAdD3VAq4CvYF0k5W7kQQdyvsyXXW6s4ExfZAdbBkoQF1eR
viAj/D+Iptr+x+WNepW+GZPit+5+tfOgABdpwIfYID6Xz09NYsl812e7KgtnCPJj3CMBKnL1dN9b
RKmnf0CtBKCwGaaP5/vpULQhKhfD9wzqHdqGggJKLoeCBJEkmKGDysY2dhNHZjo2smkBMk6lP9Js
NyzHa/OEDiyhVbWU48VuK2P5a6vuZ8INTqa4o5KW2qfMxklOeqhyyj+F8KnL7aGXCgXS9cRK0kcr
APcvue39Iuxs8Z5aKpNEQhdrAWTzBjBBYv7fEw98gLTukuUkMGZ8mAYzvpXe4X5wGZ5PvDg6OD9c
vT03KPwLtajMwe2jT/eDI1fq6IlHL2Cxoj1rZwtkdeUaC1mfNxYltQ1DGZR7f4lyxar3NHTvr/5R
k9CTOS3qQTlUgS83P7inrodrUD7F27PszZ0qV1lPuVZAsTAYRf2uWm8Y9CxPtYHBDMXyGTa0ddPJ
l0sVeNoB07qF9FbhwOsQczgQTIVdTV5/VIXAiavOC3Nlj1e6J3uiYplU6dyyVenMjqJT5JI4oRr9
O4wXbm0MZFVJDn+7A8EqkuRhNfpOQmlFRx5zRIR78gn9JCNfSkBoc68y/5P19UAo2ORNzPJdRXSA
pz72JSRKL6mDmCwyIOmcBEfAnI0aV8Is9evPE9cDr7rzgCSao/3YYUIl5JdAN4l/csE1KJce81vl
sEfEgj/Zb0/jpI2QGRo9hVaLBLcQ4xF9XL8H+BFT0tWbWJFXwQI/wdoTLwH2/oY4lAbERfwlT4J6
scBs8m+wKSAxgByG8bWJQBtDvkjFJY8KPxZWogiu/5XEdtMkb7kaMEQHz3T0LZe/cI5Z0gcuGFH/
yVTVXXQnBjqiqNvIbwYk4jrTgvGIolTfj7g+r0eMk9KaSOAxCgfNsLhyLP5q4Y5EucmYj3YOJs/X
1WSjX2jaMGw0Jy/Yns9CPxCy8Vha6XgLOAMiieVxtUGJK/Ghb35/iM07UgFN36VIR2xqQe7wrIZe
dFmNrA2aST3O8koJBqLIVy0B53SBKdOU9PXbgfswkmC168U54O2CmDF9nsIOQ4SgQlFG2Y/Q5TzX
FwsHk11jp+6L0I4qjiGM3jTjFOcVNbs66/Zkkm2jRL7et13f9jGyaaTyVQ1e7WtCa/w1hYeaqrGW
qgJJ+VXELnV4G4ie9ARKVKLljRLXIhWcTlTO7ZrUA9QwRU6jHuDZ2NKoBs1m0hBxEO6e6xS+SS8i
UOmBdH/ZQu2xI1IZzRsmbxpm9huiB+++CUFnfO7WAR5sF52EeQaCYqokYC2eL3tjVJW89k2ZvRLx
dFMbI6u7glpjgRyy4Nkdh4JALCraJ6p7y/g8diUS9ZeV2hkn4dffXDvvMJMJQwaeNj2jMJH8NtK8
PeUvAUDq2suLgv7JUN3n2EQVLhNxZK6cm4CzvqNx0Tc2kyIsC7O+eeJVinAlxMq4MZ0emK425SZ7
B3UBxKCo+7tckMN4RnKuHdSz8I11Ba9emfZSZOUYv9Otsl15g7RndBTqHm5oDLvSraXq01YpK+ni
LdQa32TYZEWhNakgUSBjXoYilpTQAyWnAW0XuEGLMs24r76T+b99CCC5oMVskbCvNcXK3YpAGTox
2/OtyjVZhNnjwss1AmnF+RMkq72qe1xy1MZlBpk/WmpZzR+3fxy8P5cbeXWZq/LV2hi60/A19fdo
h5M8b1pvOWPb1GkiRUtIm0mjtEFHvyEFgJ36MaMPd3lJt/Fj8eBkCJSHZjgzmuXK3QMlwlcmjHl1
aKNaNrHRV4kXP0np6c08MOwKxD0GwL2ZMI/n76ySUf/qc30ZJl8wBCVfMJ9EMuvXmFx9Erz8X6iO
QY3g5LRsHnUANdFfJ6zd9SJafsAtR+St8lkUnxJtyYEKYVT4BcLfvgI4PKm8RMctEZ9t0wb/l9yP
3v3uOOrJcT2LO2gVb7FhEtql5DbHLnacH0tBk9kDBuDTrhuCnNYYDb/04GJ/RjvWQcEB1cLqi8Pa
Uyzy7ntSyjwRsUb5IAZaraxjLlb3ZxCPaXMnwsEvTQztWOLiwfiapCMheThniTO1AWsV1GvIS8Xt
87+WqoJnywdI/JsnxEjE9wgR95mXbi4pXwEqv9wQUsarPxrRtqhi+7T/ndgQ+/NZO0AJArqf/qsQ
g5PU9evClDSF24l5YjY4iaLjkFVCsVQqOJYwBGm0xHXKytElKhr9Nhst62IdMJASdb4E/6e8gr+4
d0/YYLGW5dJay4P/JNtti9cvzfON1bhKGbrHH3m36Ye1Bo+tntczYfUcoCGS+u5oXfvbm1koZyyk
T5hVkTymxwcq69/sFXvBO6f253S8dZgoHVSQQB5cgjBKNof1n6wUGfBD5BiSmwoDbDohkXmjn7ha
PTdUWj4fa1g8ebqsoe26JZW9CfhAIVROTimNJBAcDlFnJhEy8rZwdVJsJimYBysUUev+dkex0CWO
l5rL29VXmysiX+HpSu1MVDoB/um+EytMd/KaTm9IoiutZiFb4rCjQFUPKWigcbdG9NbM58LueYwu
PoACInbKi89nzxJzbwWuUhelQKZnBRw2AbmLeQItpM9Xod1S7JS3hRnJGwMRpjWiMH1+kMAuHzAW
P17cYggGqVcBA5iUX9gP+mmR2hgilc7HCWqXfeIiqug/pogyVLdQIqXqCURJvfMkNkIskW96h7Of
OF413V5HsOHdvorPsW3pnfBY1LA78Olfmd5EjKwFO2z3D/Q+CbB78rE2ZbGSyKp+HKmVprb0J09S
KRgx+Og3fXeYheRj0WCsisDoballFJJKE1XVsSL5gZM5inHiIkR3qopeGpPZy915FWuGHiw6P6po
xhR2qXogOYwjaVXUxSPbDoskWD2oQpQvHyFxSvD/u32EYWC+Kf5qJaBeY6awAda4HdOdT7giEknu
3vufurHEh/28yfFUqE0e2XkQVEi81mVStpAtU6tpfJwq7Zsq5kHedIAhpHBF2VmyyzPDZoH6f3cl
W7YZKKncMBytx+J6O6R4GE0fAM0+2DcSmy4yFp7LhutfNqk29OeuZq41ntK1ENW+9EhRSA5TOO07
7JriJfE+iuvRenJQOh6suGec+L7z0pPIlw2YtDCNeE3eIzPXyXYv80s9uw8KfjL4jcLhU6tagis/
dLayYkMafp5pxazzUsfxXgAZUy8V4098Ot29F5ggcc+8dC6RKUNJ/4KC+ij7OjGc1i/am2d4Bvxz
UrgDmIdie0yoJGNGO/IXr5ndOt4QJKDeOHjhweK5jqGNEPEE8/pgVa6i0VAuresJhv5HuDto/Prd
qhG9K9LgrwI3xH4qX2Ieme0TAmMnublp0VZDk2dpKqoxQsCE8kaDiEFm69sRJfoLvO7boEwi2COI
AZp94QJuroLL76IFrqEtaLqCchSlhZiShGV/gxhdXBGnVnQxv8iBAqP4AYHSTXwpsvmhGPL1+j8A
Qa9Q1xU7g5yTPbc4PbP/7yaw+2Ww4IfKq4tKB9WHHX4DTmP0jTilkObg88eG8yuOZug1kIrJmeS9
S4nyq8xL8/fxTcQqFjT3gM0Kv3JfF0/aKzIjZQ745aHqnP0pRO8+Q20v11pWh/akPD7lHQl9trzX
pgqMGRfoKC71ax5lZ09EvtWqUvxtahYZ1mZU68jl/bvnkM3/tjk1WA0hstgIXdig1M7+/5zxTbio
jMKB6TVQluQP0GLJ+tQQPn7iOgxnzgmUtnhQIawtJcZpDjFMhBC3C1zck4H3+NqKKjRKDfLEV3dV
oMliLEYtzvtEMhgTZfbIenT41lZXKP7Fp7OFt4yQatx6Kj12oHO386ac1/b1ttTX7mb2HEE+iREJ
oh23RuV0eyu8m7Zn26IBnD+3LeNhCCI23gS9g9OlzUvF8JzgoQC9VYp7MmmUvC50nC3HpSPp+6pZ
yxjuQ/F+D0w/6OoRz3n3w1RNTXgkDd/BW6cMIRzXEXwiYBp5ROhuWTrlXdLanezfDwKEI7B9A2vR
NHBDlppP8fDGNw4yaWwqF7JwkNkxeGiZ1CAXlMfKVltLgNFmG4hhC2I6UyP2MKvvIcRkMyrd9OXY
ZeeTr8cY/l7WOxV1d1J1/7op0QJ+/Y5xdD+m8TvKEeKAfbRSq7q5HFGKuoR8gVRF1iS80lCmZ7t0
BpTfYeEhPsdGd6gAGSEuYDUWcMeEHqKbN3710xOrWFuDXEQNSRj8o6plNs4UVuCtfFRlzhiG6I8T
6hG3OGGPPV9IKN2qjl0l0o/DxyFMrZYJQJdNoNB1C8rH/xUUyuyrtSNPmwJUGGoftPIihvqsF4+e
Sq4gga4oIhhsI0sVe5m8v/KrCGQ7phvNm5B2i4dqwjZ5JIzUgwzghZPag4Eg00BdSCJO1CSJE9F+
M2H4tgcUxRDYg3xignIm4zqdc6idQO//pEr+6bTaicsb8e+VanZ8GlBTApVFt/NgfOon47jtjKsj
6LVj6fVqtaiwSxXtuDC4ydQqhYz9xM7x1NhsYHVhuweqsCrrq+w1EJK9LkLDhqHBJpOdSOZiU8Of
/u0yO5Rgo9GRBr3On/YACUeIRD1lfPT0+G73d7b/RBwOEzgmMEwEdJ4xmwi+smwJje0hwJwaeqtR
85BRFW/whDtNnTJEWDvMNEwzUp5utA4R93bebkVL3lI+zHh3aEiPcTG2rdf2+/d6NZoruS54Uk5v
zSWK6gXq1lSGaPKN2uGWMz59FDwiBuVEFhxzAknMhvZQIJ1Pq7eDlgZFYg62aorvHxxHBfYbhr5l
vJBsCzw/iLhV7R3RaHRpDzsmpJamRVZ87Udy2lqpYiqje40j3HgbIZX04OlSoe8K9Cbsjwj5tL98
FenodK2+RMKSXI5bpamHC73NmK+QCVLy49Ys5cWTHLnZ+ZVDEbjn28rAT1v4Rzl2vMr0FOT/JT3F
Qm+h3XKECurH0KnX6TUn1hpgqpUaJjoH3hRYaZID9s6znSm+B4WMfIAhFaaADQzv1SeTxfirIqCC
KW7LUEgc4hBANtBP5IQilx9eWhranurFVNvXTcvB172OXT1RC6s+W9W+U5eijcTheJGHd1M+jnpR
V9SV94HVBV/cNU7x0aCCXAYRV3gnP9TQs18gvrKZ12B8sNiHYiNWMwSkgtcwRvqANXi9iUrYR+vo
aaboduIyk2lMCE0iSF7WacESc/4rbqVwUQrHEQbE3XAO8dxDWptGjZTqxsB7VUEuG2oN0jMbnRAj
cTvKIfOYftOHnzfQdttlM28WCKoC2Aj1o6SwRHWRPD1f5HbZfo5gcssFpEAL4QDI/9MxRvVhBq4/
aHesSUVtuvJ8Zf4p0koWpIEGLMSr6meK4JAfAFq2ENxmvFXvvzAftkn7xO2vLw6FlBPAs6ODTYJ/
inYaP3rn1aeq713lWtASNBm6HGRLZSBKpSwbPzZ+Tb5eHLQk5uca4MgUdN26BWlZ++aLV4UC/Fmf
We12EjpmkWCvZiVPnHBe1qbRsbCz6ITL53ehlOiAngKtm9GkFdoUn4G4UOOJbqUXbPpdZYJmoE7r
zH9l1qkrdMTXeUgUUtru31GjFjZsum1REjqsafsGurGRiM//L2eP5WtFemcM5bzYyIo7RvuH7rgk
gwu6IH2+79sKjFsj+Es68k365x63zFvIS6rfEiieEqLowAy0/6aoOz+jJhYUAjkNQMmCtdTuy2gP
q+eIoE30ovBXpzE4YFUmrzVaSprOLeF1klolH7z1Mj0mBwh15QXy3BnOzUd0nRk9/NyinD/vURJj
CENckuTM9F1UYSekIl6V221PTT9OpPnFDDVq7id1UwWrO9P6ix+JoN66fB9pF5h/5HZCtqinM6f1
57Q4ZUjA1t0Q1iWjq3Yr26Kby3BuCAnDEVDMlCoAtnsri2EE2pvnJYPQd26bVoNk8TaGOeDSN3O/
gqEvov6AO/7Ocu4gLmTW9xpwqeytBeZtht4ubwcdOHGwmN1LdM/PSKRf8j+pEbnoXtUITw3nKR2l
QlUknOP8OYZ0XkyDJen41bc0DjGNi+BthMhdWVa9b9rEMJgPnYDppdfLmuVBNhDwXViXO1MWQyXQ
Sz3WmGOUCbOEQ1sdvlVXWEAFetWvkU7A7P9KSPj901rLpz/rShvjAfOj41NXPtmyaYTDR6lkslEQ
/Z7Hny2MSFbtgOdJBXo9ZOH9MByOYbgqos92eBA4HzipGyl5CQMuCbTh3i7UFRkhKi3K0ZY+Mv5x
uB5ByyjBx28PRcEsplSxIYwP3T9z2tYwOx/uFYrXmX1C5MvFQHFBjYHoWHO/w6rOgH8xW2fToG86
XmIYGCu1N/ECirUtSU1M0rCkTyAq6hEgPLWdYYhSsMEhLTJGr54vYdYYW02JA6BECYiflP4sS6TX
rjUf9eQESEu8tnt9GXDUJ4TvyuLD2z+GdLTH6iwscxQi1vMLwTwtA50V4ynJFLj9e3Wic2ssYYdm
BLz2C6kX04kornSRRoPM8g3Kb7axmdZdZziO+sdm+Q/jsnUP5bmab+b0/2ZIRQW5UCd+rXjnugOt
ObkxX57YtwP3AMi7DfwCjPVTIV5f/dGPy0agAkaGvwirWyQ/CHLBmZXhvcRNSbnsfuQ8XM+QH4sW
CMikYzJoghwKjm1OaJrgINuSLy9JNEahsStUCe3adXCM96wsZIuG4Q7kNGnWrINxdsE9GruGwnGR
1B1KxH+9aw2+dBm9gy4VtqBTrNjczFwk96g7MAXdRZInxIBcyX4Kwj2D3NiEa9r2a2zLIXtcgjiX
AoXJq8S5+RgLTi6xxWwK7gMGBLikwU5r6KzTQi++QlvSztyObsa5yBi7W4C/FdAMbyPLwDa3CXlT
kW9uAZWDCpFJhqzDPP3fWJbLCRDf8weqEPeMX/Cm2wJ5nKFjpXEKV/z4cJgLX9q4YrQzsBsGnt71
GF9hJbiGU8dSbofA1wwoDU7o5jBt/QMiQWTwNAtIARIX1L1cSThBHbPGECpK1uWOHKMIq4pe8KST
YxGrlWQI6/8Jrmspx2K5ykD2/GDSQELDPRPU2NsyEavHW+V5eALZMnM5MiirgeVV3XitJDn8dRM3
f3rP14ukCCwTUvHx7tdbkSVEJ5Ip3EF32qVq3nN8aeWUFS7ivOe4cG2OHpB3UTFHqBeBouBxzqFq
QJ4y1u+2+gyYXX9iR1Cc4PaFyhdn4q35yvalyZs74ozv+UNWhQTqxveQJGz7gzxH2ZKmsn4u5njp
38gQcYAeX2JvhNbtHlTG+tUlc0BP8z/AJs9TnW4/FetctYWgXpvMY1Wid+/h4rH/64BX4DKCq6Nm
CEm9gRORdGQ6nOkGxca/AetTQ/eP82pdwW2BG9XrvqUKgzFx4O0CGhWqB5cuAD7jkhac20fQhYex
ywMdyujd2wy5iAVcC50NZP+rhDEslEM1Wl352vTcKFR0APvBZv0KSpyTvn2SuusEeSWjgI+jo6NB
vDRktWO/jLkp8lr68KNvRvO2HnKWykWnEuFDi3FaZsaztgh+VzsPshir+Wra3zz/i1FZ/yBZX4+2
NsgF9xES3d+2W3DhCLwbUGrqMNQLsjyGdEo2WFyQYsmRXPX2bUiavesVGlN1Z5H9+MFnWVc5JZrD
kWcl7G+OgycI53PYZs5LFINgSW38TIwoC39Q8Qdu7vxP/ECIkxB5BE8xQyPMRbBTfyHhUCUr1thB
bqlXRKeb8OTvJ0LUUzNpDrh2QzPmGDGJVHP1iMlnCRO2vw5IJRvuZ8Asj85xjoVR/PrYNdizo6YH
a1tmqeLX3+0tuwCNIoqbpxe5/LbGlPzCTLXF36n5SnGvtkw213qigaVS42ukBvNAn2a46v0C5xNU
m8MoPC8B2Bxv5IzJWtNpu4m+qbCimkcoNIXgEhP15adbNBaBiInq/15pesoeu8dw5QJsYUnwaEro
NUA09FPkvjca+tm3J18UaTWgJX1YoSM3Yo+K4D2bakqHVrwcjBzLI1mnYvga+Y7ukLXrXFxuEo+/
JJW3YmHtQSIrnsN9iXrsYASShAziZsIlwO4Bal1VPVkobJl1JZhl1Jx2soffhxN5LcSBevQfW5Mf
ZXNzuzSmJBcKDYZcre3V4zP3A//9R35zxMbxxgAHt20Z8dCnCLZxTeONqz5n3oPgxpfnbj5LtHpi
9CNfpQb1JlINmNK1tcRtW8AUhqDPqaZwCkYbJK8GDuTK7yx+oW+nPR8VFfXosmVLSh1UYZdN3Ma4
1KgBXdDyWDXS2H1pnKfepQDYeldz2Y+5SHrHiSqiQtH+1VaCyOJI/lsbOBFuTZVfF/640OgCIBJR
MVRUe9WmV8QokdBRI+esykRsLYT8d1+bdoRMJDuuzHz5au2UKV7FF+SGtXzVFnDESDk1hV2GA6sU
QDYEeQ3Xd2qNcClnrhsIytXP0TccBZZeBNbjzhAtWbV6A3n+BKaiCXLo2Tbz62DVPmn01xshX/im
QYaem5WK8JvI5CB/2vYAhLtWcAf0w0U78+A087nGc8MI80LPfNiiK1VSmUS2q4jCHxMSIgS++LlU
pINNGwdaxrfvFunJ0hjyOK8iHAJFZG4QiOjV+M16QPSsxYn0Sbn0RwvqG63PXoIEbziHoCoshoT+
9Xg3DYw0fUU8y0sZsL4SyagohdZx5HoioGR1uqz3dGKUSU8CFWNw+OuVDxA8hZ55iCqvyPcywlaJ
/vByWnyjT9LWSV39urEkUM2wSnnG+EKDo7ZjHpcZn3vYzMaGnnfWuYBnr1SA8W0lz/+s9RzQXGQc
CjWgD0d3San0peVSPosaMHawC87z7xb3TNJ7asF+OAd2u+1EJZoVsUeWTn7C674sjclfiQo4T+z0
I9L1GCyLHMogDhMblPnw07ryZR7EDGj9BnQUz6f9D211iGM4X4NgKfM3vy80SdtAYWSOcy0kFLFk
YStdzF62bERjv11ClOFLzdb8rpH58UEI3wQqt7LUPTYsIK6fCxgXZaQh5hgNOacw5hfp4GJcEm5E
AfW7Vr+wxMgFF9YQtCJo+AKWJi8UkjXB8owJv5H5/fbCG5xkj9npvhavCNjAciWnFAd00r41n5RV
+VTldcOHRFRAdRucCV8nJ6ZYBNrWrqjAE+csvS5Ziglup32n4num+MHxwZ2vnTw1/JX78kAj1D9n
FBML1owCvqfGCp1dd5/ejfHSh/5EMeNw8s8d4E6O3XHYc5Ri7nn4c1VEd7djioQvdzWgVlduJjmW
BBdNTcP3f3Lr/lzFZiQ0LfausYtWypQs6iRCWgMVuX8L7/JGgzNBd8fkFt6E2rMWZQMwGy5R90yi
VtQldQxIINoTN2ncOEiGm4O25PXAwm0MAKjLO7FSCkgNTZ50hKPY0FpoZ/CUgxgsuRz7jQWTOaT2
BYk+gpMqCno/s6tJU3UzuG5dD+DIilKaChhZQYHIpPEkg5+wAlIvU0LFqBCjchHWKVOI6nXEEFW2
I7E4z23TOtfGlmuiPd9532L5+D0ikGCcfP6by0PxhiQtNkgkljIfyMUxw/3iCMlpPwfSE1qHpNow
hY9inLzry1FnMNo9SFgrde1mH13ahm1LTAz+bTFPaiCSjDWGMpYaGa9r1KnOf6uYIDoBjmoFJb+Q
g2LTAYX8aVivSitJ1RmNHcgEjk7SbZhsducQk/LfBKl2Vhff1mYRgGUPx0qHeppo5kGSUOgxPLzD
lvia6TRHE3/ynv5A99+wfJX+3I1fu05Tq7qBLVePCavC1CoottVV9RwWFNrIu62LPGNj9yvycDp2
aM6aubighRUaDGZcbWcQK6bLYiA83CrLUvIWsNwv4XDV3QZctdhh/8Dop9fL8E+u8P28+3zokGuD
/mPftpwMBDIdujobMrKwn7YZFrWGg+jsKPrBXON90zCSZmU4Qg7GoQJg0efFVnr0kWdTc0NF4BrO
35/DNxI/nlyC19Kyg25rU0IQkFLwvpVSOvzjdITA3scau4CN2WleUcy6FAMJxJgwlKrw8ybSVGV+
B7Qi48Ep6TqKJJcddWNgEGt2IIO1CqzjZ0HtqKDYXt7yLkXajVFx2rnwsJtrayOGY3imRTd6Gre/
zjdHFm2ShJ2Q/MxxjOcDppuFAJSeREIjOccwv3AqxmcXQQOnr4IMzfOxjN9FOCTsLbTUwlyBDECT
TGhRao9NfUq17gV9G3OtqT4WyNGnyoUzBYIve+sHv/NPcUvGzltWDfdNFl0ibp0za2ycvvf4/K4L
kEUkIig6GIRTj8IQINTBFoCGzH+7BboU7+8ciqRPZ6BjxljdnIvjvVTAf65qabpUhtkT2QVJ8w/4
65IkQRzETfmbw0P1lQGlPFMvrClcvSCAKY3jabCkTbaLreq/TePNpPzdwcrIcqtWg8kMa213nEfd
w2dZao4eV9l1EmUczynL9z3U8saAkucQX2ZURQqlQAAdxJTq0+cQwvZegu3kR8OkzaBlFj4CREkZ
1X+lsegC1n3xpWUbfz2rLVhQVOZP+w1+vgrj/I91AGiLTzyEDgNcmFKT99ca4n66FQLeH0nQx2UJ
/OTo1P2CP0UNI+Gyg9Qipjd0Xd6AzvDQaBrfuab07EQf02XvOUzRw5IkTfrHF9UBTLPDsxvJ6aeR
xAeW+9J03dmzURO0dES2tlW4vg6m4TCmdLYl8brdBRWNvqrFJQD/Q1bjSqn2QauSlQrgYqPhlmIg
6GLJZOlpqizN+94iPVpeNfDvr7cGDXWdgbid6mlQPONP6koseiA0HIqjaC0CiHBEsR7bu9vHPdzR
fLup9Wag2G+Gc9vsFZjEq8HbFz41ihM86wT7R6S0s/n8GpiiK/6Gu0Cofse1DS25FiNkgOtB5cpO
bWYIvYqS9xmlyjuQdj4V1+L6awk5iDPwlo+X375MzOIuv6XkfeWk/N2+r+Bex4Weu55oq9PyqY7o
dUCqnI33Ut+yOKMX4k3+hw9yYOfAK1+d1chIzEPqlpbaVxjyUpe2f6CJzxredzkeC5vGIBfHBrYt
LYTdj3XP7ckFtSXIK24KMS0pCTrzg3dbqBVKFuVBTlH4sDui3OwGxKDuMemLsqREFddYwTZcsVfJ
YolOf0npT6r1ERCw0RnjJKHGi9/bC/3oLwXXJCmo4q+m59+ajjozrWGGRIcPIHwzKNrd82GAsWZa
mr+jiWEt5w1cKFVRX7Av3Wi5johPAb3nr3J1tcO1AhpNDgF56KiccSYx8P3Lc9iw1P5/SKBPnCFk
eFVxD70lDFLPQ5pZ6lyUTZVjbzRY8o19miF57ONmUmEK5Jn6y3r51qVCgYoHY9XYcUnW8kyMpGVm
zfAXJIgi7R0RuBk60nObcUuso5sTsPSsg9ULQP/LZq+xD3LcH6PmiBmKRofaeieAS7AGZp6uorr8
VT0Vc9U0W9M5aqTkOHQqIsckvH2WTJm8sMlfxfINRs3o9+NAmpwNvRu8NIMhwi/KnWrgW47xef+s
fRAIZe2sZryzx+LqSKVgPxwvxNgh9iRadjH8EdSpKgYfQY7yb7De8O8cdUdgzDogdCke3J8rqdZ9
H8vu2qcR72HCTS1se9Z/eGEkiH6PiUu+qpvfE0LD9wUJYLStQWZRKpAbvklQL4W44AntlqmvhiBV
WcjxwW7ezYrarhMVQ0cMaJpO7sOvQ8Fbwjo1Rol9cDOWKVK/oWz+kNpx+oxlvIkGfwhXkrN2oum1
0Pbs/35wSxIWzg2WhxeOOgzw/EOMYX/ZsSnnjWKqVX8Oth3twSChrtAfsDmUomEx+BbFdmMrcXYk
pv1IH9KwvXn5anE7KtVp7OMWT2uXa9eK2419NganBgJ7wKGwyOHqy2rHz0vUbCKKtOnY+AGhCus8
L4CdufiJtmVdYKiIoFyB2DnQXHEQ+p/SZHBSe3tyd3yDnaWAKEgqNvBaoiTJK4WRYQqk8PxY8yIY
Lkfv6t0QHwJkS4lEeE60hiFY67Gfl73uwQ9PqdLECuOyN0F/W1wnyrs+ybh2SaLJfEgdY9eeL4Ha
tN56NqTFWA6ikAtZHU6WE5ZR8UE1p+6mnVMq4mj5CLjhm0W2g9BqGsowUR4P7zivNRUx7o7MDBMb
ZA3RE1+o5kwXUM8Pi6Mo1pWdBpgiyh8+K6rwCrNNOMP/0hAupmkP+uzChlQCHYwHKrwxuhLEoHum
J2Ve6VbQg5OOEc3TjbSj8JcPx2mrrtYLSN0qcHiMfHY/0+xK7ojvl8Sf+QVrm6/UE5kX8VRg4zqr
adtneolZlgdR1UkR/SY12DlLXxcMWUuTxhw2lQfMpzRolveYKqvZfDVhynvZmwOrA3TJIDuA5FNY
YM5Tfh8iRaIMfMD9YKOImgd00ef95hNneFbE02ybyH7QfWMX49SPhawMBMyIeOavufzvRbR4VB1y
SnjocjT5VTu7ioFsxbUx073aA7kzgP5hK1nIeadYCZWeqmaNtmQW2f0aBFpSZvmrhgfRSw2zSl8f
shwDZQe1EqQdzGi3iUqb9e5FFNf+BdVCoQomnxuHX3tnyTdqxR077wmhboQHnpnnmSGwU3Fkxa+N
x14MnhA2NEWBepRrV5XPkwFhMe0i7CyQFp2j9l4yjpdHobgfth4jOIuhF/xa12nMYYmPtedJ9fMm
vTb9ABZKqMiEvksMsQyd2KuDBD3AiLQiSAP8ywz9iex/APbMIML2OcW3i/hINUVVUX7hrGyyh71E
7Q2rCv8k/tGjqVGWvhZwglxO9Re9lw6SQ8fs8HUfdYX4vuv9L+V7gJ+rdQuF6vb9QGHCnh99kzwR
66MyG5DaBtWZnYLGs0xk70aXB2/jaA2bkqtFaZB8VTOjTh3Ksz8BQpD3pxGYxNzXLYeYtJ5WA1Qi
gCO46bYKgH3ZKcsePwbPBUQB426fJwMuSc/5ATfM4mBZ2q0ZXKP8hfbDwXP/5VzHOeNHELWComUM
YBzsl2wF6Ry4pf9KVvcidIONIa0/8Lr+zQ0o5s9+F5KVxvb/nmjNNnBabs/kvvnavcDuwL8Kc0Uh
TJg37GCqg3P/h5qqGM7bT1LBXak4lbQxE/LjBjLGyEgeNrarPqegO4VkWFpC2RHD9V0lNgLSMPZ6
E8YNivMebKeD/z6PcN4kbBfXCkhPc/HexDICOTJnqTrtMlBjZSGOsYLGj76Hnbt/aAivBGMGpdbB
VSYi7zTmcozUR1AlTAVtjsDuHgIfpQJYDD2ZPHxVQKcT35ddLwIXvO94ASFywsa7b3jIm2H00fOc
XZH7VKKQZhawP01qsr50alKC8YWQC6mfR3H8+IM3lXhG/6w/qq8iTdfUnIydvnwbTlWsRIaqUGhn
qk2uR77w5bH9ZBJAkEXp6ZEabCoJApwmsNAuBaSs4etXX+rvxLAyQUbgBfEj5Bo9kSwLHGHS7Kt2
Jx6osXdzB+0etlWD6xps9wZNj+jgErjAf2Sxxc4k4LTGVgPi3sUxw2p1Eos4HzXxlO6eTXvG/Wox
6045DAjmK5eqz0bOq0RoTtMFq2w6TDIlJ3ygn3fy6QBKrrmXDc7dJrDZEsn4eiMwnZwtgNL0oSIH
z4n+ss4l2++7C7NrsDu5XJMwWG3GbTKCvuI6jgLKsR/+MSLVQGejlqRtrvbyrgadiRV6Px006hUJ
jg7RlFm+Fgl48ywDAYtDk+NJwq7dQvT8vpS4WMBjpdlHSObq/a1F0YKz+9K0BORZi5Diux7p1SvP
AtAErCZCyWMC3Epqp1a18GZs3PlcSZyeABJ3UQzkfEskByl9zquzG9DZsUbi/DAlEoV8p7pHcdiO
vBeB3e5xzpnNAXnbM954CJdWptjGbd366GDaycUGsJ+QDVZfSU9mTDjySfEPydsltwdhFdloNwcz
Ip7s2R/qV1pbudFcZU6YWqK/Fshvna5gD18+A9/zGSeXfXPbtvlTgqulnldVLgW1BEkYXt/UyQHU
iSL1v+7Y2j1JK/QCvlz5PDNw31tDsxgJmcdKxW/4jyQjdM7yBd713uZijQFy6/hXvhWtW+ngk+3J
oqnO4cMPQmAoEeeLzWhpACi+EwKS3EDezD9aWbSIGj2x0DULPD2wPbIYY0bl98PoxNd4Haiqp6hh
qKXil8DPnjTHr8d2R+g2SoIWGIenv9JmB8jo+BI8FliCkqWY8F1l1vqVBM1y1Y47AMrukylAklC9
hduvkfO5wB61V4/60zoxSHLy1IStFYXiUBjBD5mpEojpoR2+yyLVkHT1PAbMV3AlqJ1VsTTtblsp
PNCFZz8KA+Fy0IxreEAb36AklrrpDZIZ0+xI/UsPkZAAOUlER/79qPgJJYE954e2HqHalN2vJRsS
k2kSl9ygWD00mjMn2A/y2deA+DInVa2Eum8b93UWex198urqOrP2l698PZjHipwj8Cd57gXiJtKm
nLEtEmnUFeQoCD7hRSUe8q2QOaeqI8UNMwxYkdg3bP552JSyq5xdssgwDG/jwjK77TYg5m+po5O2
4ACHNC4InZOwhpIxXsAFyh7c+7K/AHJX9v9F+tucs3XuozCIrrs6g2PBowl4NZySyMS9RsknY6VA
uoKtzD4M+nnQ7TK372IkVILI66H0XSLPd0XNHLDZ/wI5MHC1znHyFB5BOq4NHfGtOwNb0meWrknX
8elKjCDEbcSZS6F2ufRB32rz1v3gnXvr5OezcZOIGyC4ZhLhEuPuSBdfI6tRcUyQ5pJoPOyMT1jf
/Ufkaz+/GUnyBG5WgOPWWwOJ+Zbi3Gxm0bA46L8ko9/WQbaxF++KGEfCUpRkpNge8eIHJHGwEMK4
OzhI8+tUsL1NG0CLfgLMm/dmIWu0oPvejbBHmYuoxnBJfHNKXdBe1wDNy4whUZlYRvBdVsaBBZiN
1jMGJu88bnMdbY3vJInrFn7uYPAowRdYzIcnUBoAIACvfe/gn7W4ngHYXVhcavvbJEJA2lcZaccS
UZ+3d89hzJjBETC2eaUarxI1vmOkRdghNQBa86lE6UJLbnvEAqh+kv0VHOe5sTlR/C217zsWjCRI
kv9VL8g/xriqQhDd20qwx0pB+3/liHjpVVVKW8hMkxTGtSE8U1Mcri/yZgvJWjc8spUzdoC+WgD0
z0wz9msV3qh8g2B5EdiGLaTtCQDSmtKqij7Ntj7QCZNbczqAtNk6DQZYkqRFoRpgPfORaHszgkom
GY0LIAVPFBx0kYN64kSgCYInqGM+8RezVmbG/mtQs89M8YgaTFk4CxweCld4S3bjbqIIq+jGDMEs
peQc0+ktRvsSl9iJljb/3hdIPhGh8jkvuDKZ6I2fXXTvE+YA2x1qbKCfSmlbpw4r0BVRlQah2d6j
C9f1/W1wRER22ls3h1gxn7HjpKJ5jJklh101vikwdCSWRvmIPqdqbo5PrYrf3q+Ir3oMIKTm0/o1
KXUN7YWS9kxu6feAoWoJh8Yv/1I/22nV8yV41fm22+rqbya01AS1ahd4XeDom0xb5xcLIuHevh0G
Px9UxIVUEz0NKSEJTDaLphYLr/ATYs7kjmFtoyZuHw/YsRwafyyG17FBR3Jqj/XYCTPlmpGOVAFC
85MDNnAJdH8/3AcOq6zTDdiVcWbvp5+p5B2a73zYE1eAiwnCF9j5swOzIK6QPQrP5lCeGmSekriB
5SfZiaMtciM8/fpEC4Myh5G851uatR8Gbb2EKj2qPXiyBdnLS+7LKBZKr33gAl/8TpPa/ip5FwHl
9o15cYFKXaneQuIzYpbarvSupXCgta8yA696B8MNWTK+5dJ/+BpuNYei2cAzUjlUZUqm6ekBLnkb
/qictDP9ewQ+9IjFjuexUHVbxP5xZK89bSUr/gKxl+qbuYIjg9/7SvzMJNue4+e7aCNCVm0hTdaW
4f/2Y3Ju4A4kGsmjpeaDhi34A2yxRqnBjN8192kdQQKlMJhvVNkzEJCYGdLxueZZJS/VS70vkSeZ
0yqmIaRMhCbwEqn48oQvfZUWuRcTIbp1TRkGLZ+f9UswxyTHvHZSxvJBVRmpUUPMbUi7hDXlHCY9
iqshofKYuecvizeU6PYsiPueeKSaRAOUbLaA7btXL+S1XqEMmBp3EuFim/VUXt4lKnInjz6EZ3R/
xcYPMwWcE9EzI+kNeOPZSat8EXwnoF9vNvjzg+mKINCMXWtTvmXTAdzKO4gUBuBaPu9lOgqRK6pt
jw1WC39O4RCveLGXcwQDZnbAhXoCjif8twqEcuLt9MBp/92VGEMXEgU8dBLrQP9nIoArtVIIo8aD
243yR3MaLIfr6mzGC1l8zNMYE0hLX+J1Mq8IpgYfB0Zj7ZXb/LB2WrAlEMkRetiEuigM9KuYGqq7
C3inNFWXQu0drrFgsw/ryT2UaYQTzKDF4ONuJHKvXcVfy5aVvpeHlXEkfCT9lAwfALN26uv9Nizd
SCDAIsoFKtG2JSs/Dt12MAU+bmX2w9hS/qaWWKnvYJFbRA4+F+AVUyHFa7tmyvR7KAW8MCozgkfZ
5ho49rCB5+CzxW3AEfkQRcTObke1ZMzebUkgkn7Z88omsFBT9ISaoaoHRZ9eV1LyZUoc0QSk8vrB
7vlPCfaFwbsQ+/oLIZIZPPUXx3s0tC9s5rBcx40dqoEbYjxQsjZnLjveFQrYyuoD9LtNK+TFaJMd
zv6jMVHJ+YaQGRG316+tfaPI/7AuxkhAb5v4ReYTfo24HWxBjIL+fsaOgNST7AAGoaqgwlD12gkA
psKJBJEJKRb2qbTcImGLlTkH183zTA3Gv1ngVOpHerdYvfiaCcZVwX3TnmY6ZHXIZowUuNcxoDDG
dVzx9miyZOmTGCGGfFvJt82lyPnDCADkFa5PUDOU8i2vQbc8nNGI1sqfir4vCO35ck3vBAb57dV0
8qlA74yp9GHzlV7Kn9PH9K57ywYLCrK4aW9wLtSKPXytq51VJgFpx4//MHnPjLCPqJSvhCaZRPZO
cd77LWZyYvb3nZGqmBB3qMBp0+D9FXTmFx+1ib0PwhKtURUClSQGkiwoUzNjBajSa/Uvt73zcDEM
eY1oaP1DdVorI3KBLKJSaD9BfZQP7LDU1muC30mVh46V3ESfykAj/4KYpOqPES7Q+3FixIsmnMcE
wNc2I94bCCg8znjYW8n1xgbqQSdo17+Kc4MROw3Sx7KNuUFylGWEhozkXgOWPjAPEdunht2s1pQ6
iUuTd49wNe9+7hczJgv0xD9SVdQKtT5EMuEM/Z8dzpIvKvZpAxgBJe0IzYtaIdXpjx4qiB+41Mx2
Q5xfEzZBVUmBJkNb+sWFVJ6dmhOxRysUrccNQ3P8prylAce+QwQk56bCbl0gD+joZvBR4Ahd3kjc
FmXjYUTSbPOkP7ul8VPtfnY9WjIzYRJMBHtonFsd0kSoVA1XML3oHcMwOgT9zYvWXxXRVgnGFrMu
d+jLDI9WC5KrJQ0nxtcOSHQEfagdHSWmEJomee42BBRkD8x77ToYfVHOWrj/zNlvtV05p6EUN0q0
/RUvDJR1Y2TOJsXrdHD+R68vm3v4tWB8z8eaoEiATNcRzT5vSCcqKd1F7RCV7kqzTksbUl62RLB4
+06nWR5YaXHHr0cKUB7H8e8UQu54YSY8J+roYVe8DBSohKlrz01pSB4iAScGOu+PCk4tnrxich7f
9lg4ZiK5LrngpqHA7lcOV8bkD/Mtc4cS2WYBPvQYO1M93J2GiIHWa6ZlJmyRHr4SzvfHmHTR3egH
MOyJoX+URhGytFlLt8N9XovufvYsuHHMJiN8oTRyemYOUvRBAjDWKTzyhkebefeP6Oosctmp/HQc
okq2aupGyStdhj0N+AQJAvgDYIVLVC0IM6sJ6PHqPlpdWniDp/mKlUcMjA6LwZ3g5/uOLErnwMIi
nH+h7Kki5MOLgtNs0Dczb7rckM9v8TxGa34PONM9JQ7vIjSQPnhTSMg3FmWIvXGdvdWjZKUv793f
Yjv4Hlp8ebHqZAfgjQaEJIWcdyw17SHIWq7yGpCKDoWCCt2xp2eUQ8XC5RhR6TGmnVqUz4F9SOuD
dl4ukNOEyq9q4Y8YFF3ggnhUqVzQJqeaSDlkzbRUQxwGY2I1gVfdJsBAJiQY5v6Edm3YcqJijc0r
2krOiTA/XxOunuR2RXhIuClRShToqllTzzuDhO0BTgHGElfbouUTLx9FxDD2xAjCaxt3BZG8xVA2
/tTBJjTKeLltxDld644w4jKVZ7j4zoQPMtOwUhUP5DwE5Y1e3uwWY/ZploadYEsMr5apkc1bDUs/
W9PYoee1bHz4o/gn1sOIeJRjorXKCT5p9bSDlnbfY4Ylze7y8DWPv7aQ1udl/37LJw7CeOz15lDC
aq5OhAjpevQFgaKk3/tmdCMh5ZTYTZvdDHOHS0ZEHIBYp5JF9mtDPO6WkKsORLCUW9A/N4CVexNM
zITiIgYuCdzssCCPfDRg3Sv1AXcNCinod1BM8GCbKiT3BMz85Dd2I1763bhHk4MlyO9pewDByOL3
sJfH8nbC6GuJ4LY22VwZdCEgedLuPpjqKRsFh9mbB4Nrfh+GqPm8rbA6FOzg27Unyib2m5Q3LQhc
SuOvJlls2c5qPJeE63Kwp5HeM0emxjTO5DE6xrrBzhUw7hSX3dwcqsk4caiwE78jF7EAMwAafVnb
fq3dTNF9PWXVrVRDQ/PuM3CK8VqyUTIcq5/ouXTy6IzUEJ6IdwM15bifxRbgsVSxyiBoINm+aTf7
eJW/uWycYFIqZy8JwrQILta8PwfWQngYzvLt+7m+8NUskmULSQx04ApmeRMHDbBoM6iKOvNJDU9m
3ShbPvVlRsrQWueiEJ3+RYjrA5+Ph5hby+JW7SvNZUc00b5rvEBXvqLzS5Y7BOcKhKiTRi87Kzja
71mMgCbFfloqHHAaHkGNqEn/2x1fmdetvWtXmt6b0FHXhmV/N1fgZr6bMra8GCi4oLG6W0xBWX+b
lQmp+/sTQ+xaa9hBFyq7P1kCXT/5lxj4/gud/g1liTmHWWEgkroA89lOhreDyXCQR6zVJ61PMoVd
Q1GRStSlLNHoAkDaOSHFN1R4lcMZ/bJXRoDRzg9IX8EdbNfy2xZCPeJUqF6SBEo8VR72SvuMqUjC
EZejK3ZuxS6rZgN8SkVdWRAIe+QBpZaKZIm6uD40rFp2nU/XqsuBjGeqNDwgCfs2bld1VaPZguxU
2FNyW3iV8qtFR6QzP71qcCJJdjkufj3J6lT1NcIJIAvIMwzzR25Hcn3lLjNUCCyfzaSSXNaTSzsQ
rPgubac+UiNxfkndfil3Rn8IvQFBgGzCyYrvs5JqbXSUAHnWWDdAAt0UgihAhlgp+lccDo2DrEji
/9CEcz1jfOEsIJzwGsFdI6y/4+hCOC4pGaDjPUYLaPA4a0kppiY/am7W3EGvY/Bjc6gOOHdyQTls
en4oO/FUcIETwMDTVL83hhD9iAFKkJoih0j5Zn7ZwUZ1evDQQP39x/Hq/kd4DpRn5NfsEUZDh0XN
YPYH2Hw0wtrSSshl15Tzha+gBsjGWaeGWjtJTul45mW2kugAswTWVMcGKuPQlkPKcycM7LJfnGJT
KWj79dnGkBe5c+zFzSZ+I8aCY6Ewd97II8XHrdI8ncQzbspP9bWk4Jui7xO1oQWeHBSkwnWn4yto
tUjEpuAaQh8rwxAh4oNFJO0fLvlpxk8ZhU3r/joixK86vU8/+EfGbFme0skMnQ7FnbYMrVpd4pwn
//QGyeaeXdVbeSVP6jL3isd6RiBZrfhjuOV9zMBONMrqAA2oLc3gN0tdhgYCIp0tcSfnZHVg6a3m
YRzhYtjSZUcBznB9lWOmqAWRDqn35qTgTaLWCaSVKh6R5U8Y9Fj/ic05vey1qj7QDwMG4Mkm2ndO
t8b622VoSKs7l7GT7vtYxRR+kNMHZXUkOm1BdoEUndJpkKkkYWZ0a2xGXmpmKZmjDBiSBCMX+DaH
7jRPgIXncNBhIj7iI8FxH2yUvdnYXgEl0UrNI5wydwKVHYD2tCp3RjRgRaUJ6Pwa5jeVi4O6jzsO
/OVF7Ckyuvw2ir9NVya0fQQCYKT/DRqeXob6gs9ULy+//p/EANo+WsU+pyzvA2jrN1nQT7Oeat3Q
GckhkOI5OeY5hfacp34dSX20FaXBsUZ0eKGKH2s7RMSfoIi3FDGEOGzefNP8iZgAytrTNz3mbWR7
EgfbuRXemjxYFEerpnlJmIiQmxA60AfifXqLQnouC6mZ52M/Eb4Ur6BbQ4SdW0zyQ9x05OYj7x0f
W2x2KX3GD2YwF9qRethBtNNirxgsaHobzGqUpqGJoNWtNKgtLf6BRc6OigXSnBLHH9wPr2TQgHwL
IdTcj3B+8SKv2NHYI5qsbruajKoReoBgIzF3P2wUkWyElRelB6b0XQwmxUZOI3vYtR3mL2+oDI7q
KoiINFZl0o8iJEOs/sz53Sk51CjPI1ImaZJ7o6CTNh1kniQvVdP7fIUSdpFANsWagqQT+GaZNesm
nQcNSPQHisEeU3nzmHkBhSYmTXJAL/lifqdGreKvoUxAobrw1dLGFCoXlG5ctyd3tG5+MLI/2CJa
xtIDmbYRxzT1zHxsQSGSFggwQLQ8pES4/N2cDBsAqpKFZGdvTXmrKXNd4q+lWC5vEtwiM+Sbs+qd
1+FXF/fRg6F7C9F4423HocybfMeefouUS1+LftK+mD+sGEtiBt4Muswa2IyldM5v0cpvEybFWyWN
i1GDuFoKnZqkuT/v1/oW+zDQafBAAVKnP+420rH47NXhc40BuUe+z0pcyCWHXNin5G1WA/Q1y22E
8ypCvt1LceDF4uXrB7NE/Q7ZoE6mpDL8uHRDNKW1zB9KVNeuH/pQbzPa2EkeV0aY4fG6bEbfnlUs
UlJLstXktC8oKmjnYlhpQoHmHoH95SzT53e/tciiA20ZOdjt20ROUu6GIwKCHIy9sknADS439KwD
y4jSQ3+Ul+KuSqmeG8tDbTB3YgpXMfHyAKS4/uc448ws/aO9xSbYUB7n9c0Ot8qlLjQMI6WL/1po
nxl8pbwn6P5N+kjzSoqpE4yhxhdn02LePZXWGbNyzqPCSZM7JWB4c8eeF/9SXgnBFyX+nmr6o5Mo
lNnW1tuuIgzlArXZL3cxGtp0wnMhVg8/rlk4Cl2Da0rnfHCm1v4kbU/JYinnVPAMyhK+N6iUL4bF
sCkaTHDkl00uwuLaOAY9KkXCaTkLFyTQJZ9JmEjBeZ3glVNp9A+eD3S80NSYQlWV2VdxcggvdVOY
u0YPxbHvDCRijkVvXX3C6ws6N1wEHaOKS40bda/KYU5E1hfMhET/w2k0pLHq9jf2hgZ5LLayOe/d
5aeRbXDFmcRii0TdYonqaqonuGIU1FsWGIG4785eIa1iAtN1kwRMJ9TDdEJn6vT2RhzNXV6oP7ZF
xMCEA43yuH9Bgg3JBMuYl+f0qyu5pGy+XcKHHapUhmYJ+tfDGLzIRFXuelavYa5VANNiW2pJ1eJc
XeoVaCdGIyebw/tUGWYDjwX4KHNLmQmgtPXa6UMnwF0kvSrkWPQYzYxV+Q3DMt4noXFWFggqndKE
QjcXy5OlT65E3MVhbW0H5vq/ixktNpRWN6My+Su4VzJ3WGCpedV0C5z/peD+INYc3bmC5jxIign0
knIL8sE+5fSm0z2pv6IiUiPtFZKMA4nW4Wan8NGT3Gstva+VXd/AOLuQPC4tIErnINv+SHDrm1Zb
aQkDMW6Xauk2RjUKilYHAVUmatXO0vJGlCsXkvnjwDvegM+lcjLyu6o9aTwdz8SG4+UzGEKUdTTn
K70PKcdpKOLVEjB537akRlxhjFR7EaZTR6R4bVVACsD3KUJhMUMs5K2izAvtubb/9KDpIAqTxA86
FQAI71eJKBa1qMUfHMoR7vN3igF34EmgOE39O7xqnmLtXbMGnx/WQOlY2ltmHDDBkQLfoHDsnUWh
m/aq9m8FzJSHLn631sAziT4lMrGKcqeB9zK7BFKlnyWmHeDec/CX2/9YLOnlTWpp3iE9tq+jOKnO
ze2rZJWsxD3RG2QgfIXU9LRLf/7wfIDUlrK14R+P4P6HnJgd4in7vbXLnwDm9IllH/c4zZCN9/Yt
GyON9uCjlAe1UWEz8CP2qms4DgR5qtI4djedO1uEVUO/NPxKLGpzmWFoexRJE8qhbzOZ1H752zaH
mkVk39cX9U95ic00tgmsZ9sgPVbIhMUxDMpx8oZha7KT+qHC605y2PYFKKpLi2Mmuv1xdOkVDc+H
PAYWR6jWyJhLM9M17R2Igmjb1ckQoMFIX7Tfmg7FkaMD3h5B9q0HFNEARwXj7S8+oBB56r3lwu2w
zDcEjQ8sbBwWAXxNKQoEBfFXylEx9rw/qTdC6MnjWFQdv01CaG5PeUgEPWE8qkyCCu92dFcWep2r
0tZvrhsgoSwrbWdXhS61jcWuZWQ0h5wMLdDaQjeRYc9e7HT3Pw/jwt8q2kpBH3oXUwsqntiyLzvR
vrOhn0iQOF+8cJ36kWWu9hfXlMKuZvQqo7EFb4N8dHLyH0sPArmg+rk4437w2j/Z/bGbaKiWoqRj
2ghX5GBgNli3M32gsRQofewZTSeB6UeEEzg6Rk1FrMzZt9Pd/uKgGkE36JoEzlgE2gTkBm7XQvis
9Ube0uD4nRFUzX/2vPPxSvW2J2fcMk5kA75csNHYvII/b5oH2ttqsobNBXfp4s59T/I3vAFbyp11
/rMD8xwH+Y4kk1HblSM0YZUjNpjtKtFFtoJxGhK9xeJlC8zHYh01EmPVZ7TMVSUw2MK/aaWpFE5k
I0PjT72TwiIYOiplWm2HxCUZZrj2n0eO/kWBvHZk7RCiYpkSVmiCmqTTVZXP+TszSh5i6bBptrOQ
l2MkccnSF0QLTzSRm2ArmDqBUBNNSeofTnEswurZJXIcVt98KMd2UNTQMZB6Ig/UG4s4hFF/HcAy
F7VtA4+s23KPolL4nY5YxoRP5dzVelCUIa//Hyh/lHLHrIPk/m1wHHnNC/B+c1VmgZytgtmaTW5T
0VEDdiQx0LjFXb7Y9oD4cM+PiTKsXvfrLUdbPbigTaCj5MtVwpj6DG2mc3Sg3r5lsKUXB1qhMwm6
9CF/7/qcTkEwZ8QDBF5ykqw9qrRSHl9CZE2fcVNSBKp74y9LfkCyWRt84U2P5J2FcSIHzZwtNGLi
zgjmz6u2cs0vKr7HwQgjV9J1rh5+Rq2OqVUJzyveKH4kkqkWku8A0H5teUYqEkZ7FO6Texzg8Sl6
Rg2Hqaz4MsQMJre9WwXP2W40jCh9ucUVqgpstJZGhEu8+ZnG6oIrb3MsFyg2ajtTfdT1LaONE7Em
RriqbCq660Ye5gHq1+JJDFteIYEUYKprEtQncCh3R4AQJtT8KG+PWaqtd/WsLPHj8NflcV3rNY35
+6SlOPzQHuuQAAwlJcc8DZLaWe8HYiI++MrWJqoxiO7GH8Y+Iy7sjBGRx5x8ESWMneAAKrQdaq0b
FKMFkjc/65AGkIgF5fboondRhda5WmFI9V3s0cS/RhuNHj1aRCNRnhtmpMszmT6URTwTOF9TqDZ/
47tDXQVpgZ8ILyBmr2fBWHR7Oz0ipTTXG1SK3DqUMsKml8jKTvWmNIncnsylLJeLponp+EfS4bGf
CUwIL4bqu4l2VxULZujvAiRUkzS6XE1/aqZubF8c1EOfijqN7RXXyDl70lTK7oihLiLay/G4fp8D
zHoPzbH6W+IEIjFoBiMjmnEBakieO8MUJurAEW07EO3Y12bpQfgqVb0w8zGNI75GRxhc+yFrHpGm
MKM0jqN2DBkuArUTvnVb7YhBdQbMAlGFxSWU2DZi1uwkvHa/3MtYOlMG0aoqZOdlVCDYzAdMScqo
dQnG4K/dGMWyDOVdD69hRJcOh8TqF/hpKnRhQ63NnDRn7kMPqLp6KD4+Ql0U+levGgwpfKKY6MnS
EIf3cGXxAde84VSAXWYdc2mSXagWc9B40S4YDvUQ2m/k2jmpl92UX6kQngiE+WlZrweKh2RCspt2
fqIy5FMyx7HN1swCjFotA4rqsw5HP9qvpX7CKPD0dJVi4udYi6PhrGgOnWwRqHjG2MZ2CvFh8gR5
4S2CedPJBnAoUSaQzRa2DhAIqYeaqUvIGL6FH7/ZU9GZQ0tn3OxtSvfIo59CyB3biE8SgccWKr9j
9qO/xwuUIE/pss4Ynic1OfZueveTq63v3RQZhu7A7W0t+m5Sb3hxNsfLDK3BIJlWTIKg1TX1B3p5
8JW/T/OBVtI7gvh0qckgV2z/CtxG3KGp4wrGpBh+zwN+RIdaWau9vLFNAoW+dHxWrAPi2ijsioXJ
wQlaFWkakET5UFP30RN7RS6rbVfyTXYGuq0pCcfbYU4Nx+Cmo5YlyB+BhGt51E9YOsEeZy/mYCau
+APtg1+NWlDeOZXdTO9irdB11gnDD2cM6NgJgorcJ4V4icpTiO26AUdsZVAqeuGePjG5inRhwq9h
UQVjL5U6Qd5XlFIiFvs36//peiqaVPZAhiQsMgP/4UIRO8PbyRdxqayY8sBmtn+fuv+kU9UYctL4
39S7t07nJ3t2zwc/oD0zcblCNYmrVTIJ5gNdMiHN/TvZHv4fmjHx0JNWdXnoH3el4XimcZv5T2G7
0KXpzeOOlj7Xr1KmuqfCiGVW4HVDUomu5rXOmY8UOOq5MZYQwOCWXWbY5ymvREIC+YQe2518R4sA
s6UGGtIV2rbAvZe57YyAhp9rBISuHgZHuxoJftQPdNY4MkPAq46TJgDNDrz6PssgNAGsZvTPROwg
sSlCTMS+JTKE1Ykh8GWZjXj04NvNSyBt9Eh4i0xMdolXGHXKPTMMn/znuM+U8sDz0oUu+ja6LDY6
YtEOpYuev8331NG5UOisexD8YaznjFm+O5AM8y2noPmRpDHluBHRoCD0RKvGmcnqFLyFXrxWbwSz
Wf8Q+ylDTcCjIYNMZOmWUFJ4+5olQkRKTVBMiGElijvWaQltedQ8HUXIub0X0xowaVdw8lhfU+BR
SEYxIphrHCr1cTz+Yf5dEVaqzeKbKlpDHjlFgZ3xLah7+YHvc100ki0L4lK2QMbml3sDW04d5Vxj
nL06wXzxiX5oNn8uOYtIfGNqMELOMvJk1qxJWSKtERB6OeUqbgWCdkUo3k1Tg3jTZswGfSw+aBFo
SLYyqb1m8Ze2kSzd22CG00zzoGseyPhfdMHLkZ9rUf5uSkF+52ngZCLpHeJBSuMnRMNrr+bt9U2f
bZa0CgwUpfSl5IIpl9uj+lYa85OLTms0bRkI5Ojq1bucYGIqH2cbXWCUDIrK5PtoxFfmD8kGUYW3
Y0rMxIL5C78Qrqi5GyH+rOvNyxewT3zBDvFhJZ4eQ6o6l8Az/WzOy4/kUNVPCMCzkSNnvclM7d6b
9MlyDrgwmUpl1YoQNDLlVh0BEoNDLtgzUP5GCDVQGQf+TH8RC/JumU2Gh9pnPVrKQYOxV6eIcuu/
RWy4qTIHiRuzZd9yJz1VK7xq4N2poQiqD0FnPTHZbnLag+Op/XLKkmlM8IaTaLQKyAqLie5rhTfY
gdUGRGhAowM/N9ANQAsPUj/DLBMhf96dIX3IVkLjJIqq7WQg/IbXd1uHHI1PlfzN70MWiYOODn6Z
inF88zJWGP7xJpyXKwk7qJKkw70sRpYxA8HLRaQGHjndWqoTlY8oBSEMu1xLprI4F37A/1x+76Hu
NcIm7mt6LHWMkTLDr15S4c/abi0MXrkPfcs8EkeUDOJCR2GSbsLNErEyolP1OYET4sai68d2C5/B
DNOvu+DQIuR6nzXncgz1hqIxVAWoRJCCOhGlfPWsLd+BtaG/BSeEd/IEd+ZdSPFmm+N0mhZZ08LU
FAQcgYvidhM+3oefiH+Fenv/SwbQmGskOa6qDQb5/CpeRLUa5joWQd+dQZtFHFOtrmxVBua8Q8B6
Zo1T/PPTnVwrbRA97DIaXEFKx32yIxwp9l7oI3W5OgfaOlpdYfmN+TCwT/u+aUa0Rm9c3lUVSPvz
mCj49W4PbP3rl4QAhdkJ0uZQdNY2/DE2FiFuCUZ/m9zTpMqzOZBulFDnrV76sZ/dJiG3BxTSJ3Wb
ckbA9v5d8QJj2sTAtLyh+bJvG9z0Mt74V5MYEjlcEhSPH1pfMbjSisomtSTID5o69d3ggK27prxd
HMOd4LBCwVQPvsWoujhf0UMIS8J4aNVKHmRqxEEFqEG0ZeV6W54xyAlrn9O1FmsxFpvmglsP4tFr
XS3hupamboVH2ohKiyFmBHhha0Xt/yRhn/8xYe1FlqPwrasvQRo7sX9myYjmWAEJ1Xb3Za+KX5st
s6pW3MIHkV6OQ2GblcRJRwwXIiki8QiBdUyzI/kiHR0d/RrcNxL6B9KHWDg7gAgAX6rlLEpS6iai
tNcoTiLMHRvz69QGCSKUhIS/weVqsvXZUZMtAeIgOap7JfiVX4gNOfEyxIp1BCFF0RcJTA7cJYAm
9AZIJhpKIky/ckUlamj8bRN99RPlHwXBY9BQ+l0zy1SzNjEN0ihi010jejOynGFJXZyQIJGMcEWy
Dzvt61NoMpkhhiOzZgRw2JIOBViFQT9O3UMg8+WS7Bqz45WzUi7rEmDBM/Q35bCDf/PSF1UlwKTL
LDNG8vkluXsHqrFnu/EpAtbH3u5ehVDNK1tVd0cjsi/tZ5LGkxbhz61jqfVvzLYf++1VLMm+mfj6
HfDvWtydRqGvuLTx0KNjv/ne5ET5DrhhHKttS+g1uDXiHVEVXBCabVODs0czS82EvZHy/z2d/csY
j6oxrnyBbU76k74d0AgxnTzaMTSBWqfeZKMNn6a/rQodK3+rDT1n40Z5BpJl5dwadFpAW04/+VTL
gbevoAr7zj6zXFjmkrY+OpRb5BXyDE+gHKeQz+4AazU+Sh8hTGjm5J0P8Y2t9+j8KW/ZZfxQvjS1
rvAmyrX5Vm8wQjfIZ7LI+nih1aRms42nHuWIjRqxBQyvQNA01VaYopDX0Ro0z5lwz8uZ9CKFB/D/
lrCg21KDcrTgSF789Zk79aCyJ2c/fS/UQbag8yOMAzf/QuuLiObp/UyFlcDsVenT507Ui34AkfN6
2BJoH4SghE8HcTo6Khh3vR+FfHe2JpwNgpP1HiORYofLAAp5JKusG5sWcPYVEhduwxLDNoVSaI+D
/+b+ePVoZx4h5U8h1jKhzS8ydXnR3IGrfXTRszhUjhPsN0CCG6Q0bHLltVXfCQ5UEnRbUu6oSKK3
YSTnKBj4AuMkvg3T2SoarSVekJ6lA0L75GXhJFpohtvnG6QvI+2GWJzmNEczxwkM3ZBsc/jKYqM1
vDIVRp0wZsO4bjGtkzRJRhiQxA/WOFNKDCtT2szMQH1/NE5C1mr9YM4yF6hYKJ5HJVD54RTco+im
XJsOqEzesWzsFkSno9Kb/U/WLyNFGmLSqHc6pW4AgqxCss+CSUVSd9G+pzjJ3Ttit/6vrYoeX0EM
9BbNfTyrzIts4D514WRYGoTz4VfxppNmhC5jH6wwjFrBh0B07MjrYLoWQmnN3LWHE+f31rcJEgao
ycP7pYiB6c9kp/+X9syuwogfZlyHFMmSRqqGQ9kYtUGCiLHW4P/84Iq1tOFxx9KbpPAwImstGZuG
AfXS8Psof8omSi3ThDKuwyhGiQz2t/GxBdYPzVAJ1DYj7uX0W2Tis74Jmz1C/SQpyhnFuNVwO/s1
1wg6KvmO7Byvh+nHy9WmiYjR6EFHYseXB4mOJAiImH599YtDk6is2iEGYGkVJ+3XauZXytgy1S70
v6Uijx5S/Q+3E0lhpojEGL1NWO9j1IFryNAidocO0RPcOvWuvjAUrwO+adVfn/2NguFDJYpLy0rg
oai5wVemSMps9Ed3pTOjxTv2mPAwA0pFECJgRZihmx57UaET31KQ1yea+U2Qi7q3lXz0YitxvmRw
YDy50TblJlBcNSYS/aDE07Kh4VKzUCgn+Z71/kG/YG+1oj0MBVIupYlPF0uWruQED661IgJwojfB
9UTJ2fkigjIyTef+5y21roHABa1ZGMDrL9sm2WFcbAuEPWlcqnOUuhiaAB8vWlU1VlFMiLPC4lpm
9egm2TYnInEgl5wrp3k85LTrqExmZXRKuqVI78jbbnTRujyQpDp5/Pz6sOSdfEDsUKOLJd5SuQ5a
80xbJtj2Bjq2s5JlEXTAfXHnvxxLwBb83nSv1d+oG9SVsEk+nZlnJfeNru2FOzMP1USfPNCYqG9L
DfOkJTwG2vC17SXscRd3VTsMb4HDrAa/Y2uM2YEfmrbpMvvzPj9IU3aYwVasEIkFJB+lEpjLTche
G4KkElFLOluZTzy+gfc0Wo85qqRput2ImetHweSUmOgj1m9iCf519LGE23ky1mqS5aiTdGQc11zq
g8xJ6o3KCT+B2Z71MQePxftpEKwqMxtpcAd0OUe26S3dmHjjTRSCzArSigf/OIBYvNA2dVHiFPap
6XSrZTVJg6pXCkh1AWfZaBFV4k9I3+424eCd5HgSU19aP7dNeVAUayxE8gwwPEz7hftyffNk09Xk
cIVhl8ErpRPpkAjNtM2PFqHvTR8x133eeHdp8bpAa50IaU5KjfErwfN19l+ZyVIEfc5jcralchcz
gczS2rljlCBE6ILaECFDS2f9zmwFhlsZjwpp97XcJCr4ui4ZxgUwkVOMtedGGfZNAQdpbvSWv1Oy
4s9V/iPBtAvmuahaV9zNv0luA/4zTLtpipp3nWXqywL0rJREHG/e/zf+6qKb3zYu07v6Aec87Wck
MfxkLCYApllfYNixDWeyRxzEGAmCuMbiEzXkek+PA2FSPYh3OTtp5Cft4Ycu5ATmXOCC3FuuXOol
8+VhXVWkaPtk2JZ7qi5IdzIMFxZyhn1yc5JRuLjdEP3ziXeg26Tfow+KUI1BZd8QT2QxgCodEG2D
wxU6TkIj9IerLbXgiiqxaxecCBKojewMWrw83dljo3f2a0XlH8ROwTTaAsESzNqrfdoA7haMWWw9
DLXATHdI0MoZ6OnLgkMEeQHacPfgEN+yHFCm5v6QH0N7Wq6ZVVcZH5VDN5gxyGHTLz1u/V7+Jh4l
qDqGm7ClSuwiEG1iuVMFULp1AfjnU+UO0w7a2tVCke+kFF44fLe8gC6grEoIcFy3TMTC3RfR1WVX
veneCIr4uNXHZUKceCATDGhAEdBX/MCRfI8X4RqBAq5XRvfwdNjC23A9VTzCt8SR4aaJ4Y0YwLFx
GsQHSOY163jLF9+ZrokGVoVRb/oO3GmwyoHOlJsKCxSlU2tktWi3v8/09QoQglNENws7LCk6kuSI
NOeVW0gEV4i8skt6JBsg8Hxks87uGAqjl8t5bsP6eQZSsX5L7L2HxZBooCDD4iVlsWZ1kxHlb93k
s8o7qCki+1GFPeCQdDqYOXLBp7dwJwmWPp+C6OEgGMj93kxlSwvEFDx4OMmpyvVn1HLgHE9WwmJW
BCcUHOaaEeVszYFsMNOGIqO8z1fO1JM7ua9c3n3QBe9uAe6JPIgh5I50kNyq7WStkR317Ib1JoKk
m6Hp+i7HyJ48i+U+5nhVx/m0f9qZ6DInXrxvOXcqOyzbhIc6WKN17K5kLjaASudRj8xsi+EmndaD
toKiNUOSEiC1uY4n0diEDwV+C4i7LbP5cONeXIJbq560wUGGtRJ3blJ9xgtw7oUIfj4a2dzFhSML
z/y8Vhq+TwO9PO+6zfcMsIldOC2t65GWK2If8/k38cNlIv33lknZFfivUaA2NDczTN6C8las1kze
fwXhpOvgyAn1dA4j/buEKnTqyFZhqctCNbvV9xMSazXVlcX6LGI/ScRRLBx7vsY5AzLLcWyRos8k
8TM8/P0IbLaOZxoR0Ek8nPlIpln0ktsFAFpQvnVTLEvlaNF8Je+eVHLbE3zhGVt4WzvK1yD4RLRe
zOK4lfjhYrfnp31qvBWkveQ/fZlXmCxIo7p8o2EIMs6yw4kTHqTl2qBVstVadD/HlLc+9EqlYJjZ
/SUJPGS6z7SmGF3D67SsOL9P6phgLaPtX0myAcHs+vLhROwczWXD7dXwrxM9bvCBOuxdckx8PRXR
oF/04uMs3JCSqEp26XFF+xcY04BcnZKbrwDyICTi2WRAEXDede9E97/Ly1iMLj+kWHIq2YRc7F8F
ECWRHIO5TTs/XYlFrjqT/HDoKax/7C8zy2rDYGTusLevcZsoPtiBhGyng7TDQXjMzckVNVGm/WP0
xV7bFTFfuwYGpUdv85qGaQuVYd4NYL2W0C86pl0Go3tg7kmJQkF/FkQ/hraSNPsnxRzmouPkqD79
u9Fima7I12OcqKaCI7f/6GuZAyloMjbrTkpHQg/BeOomTLwxA5r87SVP7ktoU060sWo7Ws73FlPV
UBbmd0E5hmDizUscJVR63SkRRTEhhfa+7+eQdDBiIW/a8Q6zgmLyAEHEBjL9VjnmKeA055hCIJ1q
bMVz7v68eIanxkCdJzIxjvT/g8GULiLnxk+1mP3wf6SNRTZZgyM409Iql7O9GFtY6FloeTxMnxJF
MefMBTDq4Ih2Xb7ohtsGmY5yAag5bndJVejSeEhptGer5cPOEg17b0cOjZJCVcow3VfiU6pcihZM
plzY3NJlUYQQEqClOwAK6YFBn3u0+WH5IaPi5aMfaxJZ6CVOJpkZwJ5bfPYYOz/B99nj84HPIYrl
F45+nvrPM9BwEAk9rL28F4b30j3xITRflapcfzMgzlTCatgWmd6uIGrYqZ66N10XqEpwmRWi8gWA
uooBDj2RAkJhwDedsKLxoIQgplE1ijF82B+mepAaOOLkslYJyK0OCK+2B4OzOa+G4MwvulEPEDD8
vBQ6VRdAOr00plYPyRjWPNUyDY8Poo0p8P4TJvp8oubfItKynqhhJcDDZxpFC+xXDMmgbZz7BNPR
h/pviw27PQ6B57GsIBDotMSmtAO/rSTboCh7q8+ROwEeC16r4emtrgz+vdN6wM5KMZiDS62x6f/L
7g/pLuxddldUKf9QbLrBWcoKkGhAO75p3h/5YURZYSZK6Y05/4hEPsCf8Nv6PFGpctOEJuZHLJLU
//fLdgpFRqBErh3tbMnOni2RxzMlIUF5p1XvsSQ2wKwS0o3Yg5NfgznFc3H0mOsDK0hY0dIuhH2X
8U1CfgY6i76flLYb+xfa0Pimi6sTk2qpnHoUvArFSOpVvUmddHfXNWiT71Bshxg6PUxpT0ZDDaii
e6Vp6GZccangU+EiYFo46id79wZYcXC7tGjjy/+6kCWXYUbXr0U3qPz9Hj4daJlNoaojdle+PqED
1OOe3dA11v6lsmyquC+XFRtJFQiv8XonKZnxuyrMKWPCjn17kHpIm7uBfroXpA4VS95XCBA5IfmI
v/sIcVMtlT3azy1JuQ2uOI1R/SP74PRND7jTm0oU1rxlsa97hhfBe/P7XW0KYIfBSb6BARXT1mhF
LYhOO2jnABs0ZumqcX3NQdybsZM5EwHgfDen/98k+EQVWo1NcMoFV3BXrkRj/aewSoRIpjFar5AJ
NC9oQJJu7cDVH2mpx/ZyC+NNcJi8xJpFIjLwZQNkXoPyeghOZlKRUtBRnDP6SO7kOk/j0i9/Kwbu
9bSNIIUFKG6EpeujY8DnO581rW5wDOC9ByAkUG1vftVQnPLWmcAzm1E7P2xe3U1TKD201O2El3sA
5cX81Lrb2gMueUVbB+aThOu6Rr+JyQS6AwLkYDeFZbwWfGWYA0g8fImsbwOemcRjoOIkNZhrsVgL
rvXeS0Aa6LusACkKktt32EhOEQVv2qkY2ptQ+5U6Us02I82ur7XpvROzHzH1xm2mrOYkU9cXPlz7
iFDOUURHYC00H+bZrodMi49KaChdN1gnthPN7lxMpDFV4XrSXTYCku1vbHnJu3/dme8gWD5hl0PR
GDHU20I4kKU3myMlZa21HqVl6hM9bksXfc140JjVPhBtfnn5wAKenkHePC9I7a9Tvi451U4b0pgA
kPSste6+crecobxSOYiRibD2WiAp3TWyZigba1QQWnADA/AvqGfIMOTXmBGR6NfQQloU+3l15mDX
LCcNvNkNqE4OjAcwwsPq19T2hH1WdCINTXe9Y9rjK5zeeofx/WxZiM/dNVyPZD2yTaaeNNlNfxra
6GblXuZ0PDgbT03Xck5xAAtfAiC/f8Zmtg2BlwXGt0bvu1iluceVAEhlBIwM2qf+dI2u9VPdlJF0
FJK7Zp+m+kt+2i51jcQzG2oaZ0JjZbX+yJXymXanzvosvP+TnoyMYeW9y9Ov9OLW0ZynXfpdAU+q
NPT63/2LtiGQtruP9RJVTwPYCN0Gsve9Gx1ivm84JEgLXCVmQ1lLd1yjD3tPAZeWWHd6smuuySei
oWN76td/6ctf4lIAUTUV5wLF7j8HR/fXjxgpjY9ikezOO9Ucg8ZgsBWd5aF7MjTVB5MFmv6ePpig
XlA1v0MWf1MD9TBKW/x148QP7Nf6XQlnmlORPDHg8OG1SFfWzkAuGRCvx1eJKUsNTPtCMIpBUILs
+AW8veveeVP6vt2LuNg6LUpMYIbd+7UqtvuVvROdYshfNbMix4Jmcio3Bq96uX7AmCGBaLH3YxqK
JPpC+Cdeacxesekw8+iiN/QJ+tESIHyJaXgSeLJ7hyBeE1279rGcBZJmENchU/uGyWUqgjILJXRI
Q5L34qXk+rn3hUzIeG2wbTP1YAPa8eCKqlrdI2rxpMZwR0GzUrBH/DQTKv9U3UFwPLGB+GutPqbg
m7OWJgPhR5sX0QPufW4J6dLVaSw7+4ok5Gb5ot2z0LuXXxCOl1eiH+rWSv0UcocC/oZ1wMUdumSL
A7L5E0O+x2vqpYmEGecKP6p7kUr+HICPc8OFwSrod/EKmIrw0FGe73VcKbG6QegMQ5oL5LimnpXb
9ABr6jriAtF51Dl3nUkxMYiSXxiIAIhjuBXgUwJCECYNaceui8kgOGE8TrwmAAg/5kpNMAdGf4IT
gJe5gLuw4lWR5XdnWKSI1uSKix21LhloTiMrClxELBehq45pQ4/xOgEyU1MO3x3XBihVrEW/E6/d
HZbVYTDE5lSdYNNYqjiHC6zERVr5tCDNI0u4lTwMVNPaXCUitiVbeEj7nCFlsrxl5l1Y3Tzlcrxg
ivRzYx/T7gsw72B3o4TB7j5Z19Ghli+uefKSKRyhyA8R48b8NuRfybcdY1BTSau0NRI/BZ4RDt32
7XI4k0h51+F4E4VRf3iYzTJ1PYo/8Tg7RuB2msyABbPQny+6+hqLKXSnfi7NCInyTISiofv1dvJU
mPmMnWohJRGNC+GN9nVJtzJsoRwY9g/Q3UzXoGIsmZorq2sOy2vONOaQxaoUf4TCFU2zvkzP4nCG
uJvzGvJHodfwA3+BEbSuXUUB6uvbY060OwjHylHtmd3e7AdvasSdOdMlCjmr/pL24LjYIiQk6F+n
BRs5cirO8zHBbOxqeRUZz1NCWZUmyeXroF29qlHMN1txhRxkG4EGhG1Ayzwl/6mK3vWnEQTSTW1U
kbFrl+Tan9+dVUdzTRbXTVWBvYpn3lnDB2YMU+qxTQZ0mjj18Ndtm0UJ/puqh2/vlxJb2o/9jJDT
SAHNR2+yhb4gjf5f7ggYU88lhkmHsqKApklfeA5cTlxnTyb+jXl4ic/GfcoErqtUiLaZM4q0Uqgx
3KZ5YSvbQlJMe1G9PtQiUHIQjvWkbkR4zhfBdhhMG3ktrVi8BkLXUTb6rfBljQuCVpsSsuWQyaF/
8I1FGOxMOPkqIu0u4Qx+Kn1SB7JMry8S1eqfVfb4znr1gljPJiBN8yFz5Qoc2UqkpBSu4D+ujKDk
iAAd22rz3s/5l5ezt1RiqwclcQGAdEeSRnS9Zo0KoRnim+32hrifPkulMpN2oAm+V/jzdmsVUBv2
vugtX8izd/UcgFqoXrHE5If6ZqTuGPfbN1GaChEkTo8Ra+Abq8X9xGeduOoIEJdL0EtwMHReN/Ns
Ow9NHB5p9fMlz8G6MCR5Jx8OH0aP1XYdy1Wip8Dauvrt6jM6Pnemuxe+qp32ZUSGO+VlvRjN2FVd
E7wkuMkgFJAIddKS2t5IxWEk/kfAxYW1ubGVTT7RHoYcX/XPoTMaAPsuBbwkMfvBvm3BLrEvxiNR
dScrbGj5Idq2rgZb4k/ItT+Gq89ftsF7G5GG7/mngmZbczpe+e8sMQX9mquzoRLehnQa2PVXRrE4
6TRKjodapCupbklKH+A1S2tDnQJhc3ghIJKcSkOGqwmrXjh+inJstxp5VNg7Y4VgOYiqXdno615q
jc8n21dJVAquC4iQPLM08pPXIBxvRBfn/5HJxLYv1fB2k5ojOFE602j8sTVvEr311H9dWmmVwA9Y
XLxAXYQL5ROXCryyl6d482uqwNhxhchT4r1PIba4sPzZv1mFXFAFlMFG/KLGLLnpHy8NOvl6MG0v
HjpcAYYz84S5OesIBeSBQ1eRpD3at/tOr/qvBbGWj4lgzJZFIeQGf0CqK/Xa8Kuuugq+U2Ofzd21
mCUDqAzy14ensd7iQl9kizc6k6knosITk9rJCtE3/i6pI7BIFak2cdaN42dZQ/lBqCatzCG5DnwP
Lp027e9BnPZJpO1Rapq6k3qEikzpwZg+lJ75Zvh2nZI1R5FIOU8vcXcRwB/yUQulZFAW21oVbhYl
YeuXDGJ/r8o2Q2uwtTUsCnVegXlTgwkduY9roYcD2DtlcyMEndLLN6yFKkIwmsQW0G6n6ihq0D8Z
XqM4wnjJ0gC04msskiB70Ud1tLQcUaQ9Alkp5dngWVti+/b0tXscUXAENn8zQf+HVzBsjX2GNYhP
8RQ2G7Hu0YU5CO7v/q8Fhep9EZNoOHq4CDEfPy9IgwAAiso5HEN0t5vDlXC9f6uT7a15XZ++9qsM
JJZ/+ieD6bmeiy5WVlI+l9wkrBR+cqsC6ixNFNllgDpau5pgLbqLxV41jFCXM7J+WxP7dVJVD6sl
U1mnwKl4s7/8MxXdSBLEdvyBfvsJgNlGgt2TcY6MqqEXj8V3Ru4emqxt1S8qlcuReXzDWJyRtKdg
+birled97AN3Bvx3iNZUpEmAaSV+QhR5qdjocDgqTeZh5nHjk/bjqchFKYObhGhcdwA5o/5lIVbH
To2xDXnq1ngUf43Jo74eKAkYwNVdj6k8ySW1+9TkdJo9NdbOSw5676hTHvwy1/SgKzH4pE0Ekf3x
lEiH9ObNRPRBDVxjfQI71KEr/OUyzBtEdaClZ4XTE06oBmiv4L9f2ymNQ/8Pg21BzhC85vY89h+B
k5ZLCQQgk/FCixTnw2Iq6nIAO/+wyIb+FAHD7I/sU20l2XXksCHBDPEo4n5jYPZ24GjfxC74PgA8
lp6jW7EAibR7q5L6p1ID/+uCpGVmJCgVaCB4X8RA8haUYT+T0uRhTspFBLbwHi57/cUsjg7HG48L
F2pkjXKKhcGbnBVfkkpfL0MQihtTuTemUXWdgGjw70PLA/4NZZMhh7EhCf7vAqzh1Pa7jRqO8xL4
r1UQ5ktOGtQBBZ29HPjp7I+fzVHE9nexEPP6Ae3Snf6Xi4RJcepX37R2k3rAlIIJVx7KOvOAjED3
wc0WJT5kmgh1IpFQ0OFEN5oe0AvlHiXvffwjN6T2KdGr07ym/uz1qqBkkK97QEM7oNmY23yNSKtt
sZffKYkXSR7zogmBfQhGnlEZlKFZH1UN/rZqBrGjVv1kRzRMl0DZBQ+9bp1kuMJnb4ptp0XY1c75
cIiZvsfM5Qpur/9F6yNWu0WQ4Y3lgUdnC5Y6dIl6PPpyvXy4A7LFAzkJZyGxJxciGTxmAV1wr29S
Ue6uVf4wRdoHnch3cy/gRtEK2ASyf6L8B4R6Go/dFAE8SoJtv5jLgzUwSR6yAXWMjg5wxEFwsJaC
uvY26JSlZF2j1Gk/hv1iO4rJqiYjSskQVqqAacIU5DK8gnPLAXHs87eBGfYXK3LYm7GwD10LgyNX
S1BiL/DC/Qle6YfpyX2eTqyw/LZM0KahW+NxnZmUG2KGn04/J86C/0a/bSlwUZwsOJxxF1XjI9dr
oMxHcwV/8DyT/5ziimEYEdPyj/bePteGWzROsOrvuFT8n322ekLmNlp6TIDRzzoc/WRGmidX1GQS
JZJqdetUcrPF9kaFE9uMf2S8YcASZVBLyvjiu4/ek7CGpIsZOUVjzw60KoGpQ/ppiNnzA/Iv4Fkl
qWiA4f4rWuh6luiIqbdlHCK+3rtAZkSfRp7OcuPu667SSeoomO0/05C1UxgnBnvFjHHKx0qVgMei
SdoT5zKwLvqdf8U7AsyhJrN2QeAXENAHplv7baF1It9JB5YN3KR55LtGvFRChRdKzW2vGe6EyT7D
6u0gkIsLU6fTpnBUJltSb4nzCa0/W7LHFOfCUgFtRTWFhln/2TifW86WnN+UKbe1Vrmp4XWngnxK
S3vFr7cn/OhCfvm/SI7AIT32JYaKlHKjz9zZxQmLfYkPuXw2VCfWY8n56HfEqCGXgNQAZUZXw0pF
qW0iHXy+oyn1Yb65czf5in414AUnflEN5s7lxg5NfDnyWYynhvRkCVJIXjDeUBGElWUmuELKLHAw
6W91lE2/I68OYvVMoxIS81WY+w3BRllI9ObBdiZmUUvH9jsym1Jv2fM/ogDefTbJAolbwpk/bgMx
SZB6hYjZkSFvvczcf6+PbAPeY72j4vs3iW2mPuOTjUJ5pS+PFw/d7DNW60+EKU7sbRkeybWMPm84
OtLjE5zzWvg8KFBcUMQkX3unOLgeryiG/RgypxMrcpBoQ6+/kC2UiapiQKjr1YOFnXR10juiw8hD
4qXNFu9s3P2hornQW3B5IylUwmYt/3U7OWXXV7KLz/69I+BDK+mxkjpJW/V2RskTKBdc+AiCS6yV
VFbsmOMLdJbUyOHj/WCNTj8Tn7T3DztcU0hb2Kjd3/v4m8W5OC2TyexKKgZyH4bSKJ2UQ/grp/Pf
Aq1fNl3xSHFP7vELjYNUeD/nuJSF6SYWM9JBb2+2TeXoY1cRaFEh7QiI3fsgN9twcWqQp8uYQfBp
zgUDOjIpi4qRo7BZEsGpLHkBmjF164oeUrElf0LEEgzUHVvWF+JxUARh+PqyQl1b8XVMbRogno15
+6hJM/4yGZlgW0HZzbpgA4IKoJ8rIiZa0WikOHs36p++wdnZp5kNc/SZxs68ykRu0HtrehJ4KhqJ
+gQPNc74vpwnr9+SD8knJdvcZMI3aM1qdHjVnwf/JsU2WUIlg8LTOPe8nM9fLKWe/EdJvtpZYXV2
+v3DodZupIwM/DmwYqbr2wKTT7WHo6j1Zt5rznz2v8LK79H3o3Y/D5sCjSUybYDSKBf5wWBax22y
0QJJZfpBc1TFGooicQB1NSzUDlbBkdgTm5dxAYAczYvVfb+hv1e/+Xm8xjf6gsWMfKjW9yp9y9x9
YKYIQlmPYEW0YeH58QlTAYcqmMycv6Pa54mp2H3NEyuVDqYb5xmNNBkZjWa8V/HsMCY0dGJFR2ON
ne1G4IEtMZwkQLOeXoYsqwRIiIheuusVffNL9cxJMbAYtTNfJLt3/MsKwYltkeKPLjxgPb/0B07i
eIZ/vo3xQlhsTRqUhjh11qSQAYDWB3UoGwE6kHq0DRqnnir82t49CnmwZauqKt2GGWIEHfECKc2M
xrbHvI2jlt1Y0Ogu34PjK1Jh4/fMSGQDBY7NzAqKz8cZj9i/EvPkZOwcd61rvCkVI4vGn1xCWQaO
j22qdDtYNoreCw4A1RxHuCEQXARo2zncOEqNdm2MuwxjkptkcazJ3kW5oqfR3XQWf+UQn3T9xnj2
Z9imceroE01/1HYcK9wdCLf+Ujjv2XhjV8hauJMNzcdme1+mw60MGZe25TZWEdT0cxJKXS3aen6G
xBX8IFt2BfIug3lGuM2cj8yvJ4nXJFLIHJ9olhdr7dbExZXLOEq6qJcwQsWKPW3f92NsmPOy6JHk
259K0HwPqzpfkPGPSO05ppzdwUGNMjSiJXzhzO24EnCyBXpA/R6InLvlPrv24R3KnOn9v4fcO/8J
JMdy2wIkBGElCA8VKZtCohXmu4ZDIQJBePj+yqM78HAgHK6O2kB1OD7UJm0sUtUI+TxXq3T2WoQO
z1aB/Cv6DMyBav/VBtZQM7vqBnvimW/eSG4Z9u3s++fQdVgjmf0xn8xkQgQgGqqslGrrOL81t+V1
91SeUYIAlVIwaB2fxzKQiXU15H7Nq80UHhcbfEHk9H2f+fsmgHnk
`protect end_protected
